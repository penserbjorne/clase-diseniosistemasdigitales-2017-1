library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(10 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom;

architecture arch of rom is
    type memoria_rom is array (0 to 2047) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"800", x"806", x"80c", x"812", x"819", x"81f", x"825", x"82b",
        x"832", x"838", x"83e", x"845", x"84b", x"851", x"857", x"85e",
        x"864", x"86a", x"871", x"877", x"87d", x"883", x"88a", x"890",
        x"896", x"89c", x"8a3", x"8a9", x"8af", x"8b6", x"8bc", x"8c2",
        x"8c8", x"8cf", x"8d5", x"8db", x"8e1", x"8e8", x"8ee", x"8f4",
        x"8fa", x"900", x"907", x"90d", x"913", x"919", x"920", x"926",
        x"92c", x"932", x"939", x"93f", x"945", x"94b", x"951", x"958",
        x"95e", x"964", x"96a", x"970", x"976", x"97d", x"983", x"989",
        x"98f", x"995", x"99b", x"9a2", x"9a8", x"9ae", x"9b4", x"9ba",
        x"9c0", x"9c6", x"9cd", x"9d3", x"9d9", x"9df", x"9e5", x"9eb",
        x"9f1", x"9f7", x"9fd", x"a04", x"a0a", x"a10", x"a16", x"a1c",
        x"a22", x"a28", x"a2e", x"a34", x"a3a", x"a40", x"a46", x"a4c",
        x"a52", x"a58", x"a5e", x"a64", x"a6a", x"a70", x"a76", x"a7c",
        x"a82", x"a88", x"a8e", x"a94", x"a9a", x"aa0", x"aa6", x"aac",
        x"ab2", x"ab8", x"abd", x"ac3", x"ac9", x"acf", x"ad5", x"adb",
        x"ae1", x"ae7", x"aec", x"af2", x"af8", x"afe", x"b04", x"b0a",
        x"b0f", x"b15", x"b1b", x"b21", x"b27", x"b2c", x"b32", x"b38",
        x"b3e", x"b43", x"b49", x"b4f", x"b55", x"b5a", x"b60", x"b66",
        x"b6b", x"b71", x"b77", x"b7c", x"b82", x"b88", x"b8d", x"b93",
        x"b98", x"b9e", x"ba4", x"ba9", x"baf", x"bb4", x"bba", x"bc0",
        x"bc5", x"bcb", x"bd0", x"bd6", x"bdb", x"be1", x"be6", x"bec",
        x"bf1", x"bf7", x"bfc", x"c02", x"c07", x"c0c", x"c12", x"c17",
        x"c1d", x"c22", x"c27", x"c2d", x"c32", x"c37", x"c3d", x"c42",
        x"c47", x"c4d", x"c52", x"c57", x"c5d", x"c62", x"c67", x"c6c",
        x"c72", x"c77", x"c7c", x"c81", x"c86", x"c8c", x"c91", x"c96",
        x"c9b", x"ca0", x"ca5", x"caa", x"caf", x"cb5", x"cba", x"cbf",
        x"cc4", x"cc9", x"cce", x"cd3", x"cd8", x"cdd", x"ce2", x"ce7",
        x"cec", x"cf1", x"cf6", x"cfb", x"cff", x"d04", x"d09", x"d0e",
        x"d13", x"d18", x"d1d", x"d21", x"d26", x"d2b", x"d30", x"d35",
        x"d39", x"d3e", x"d43", x"d48", x"d4c", x"d51", x"d56", x"d5a",
        x"d5f", x"d64", x"d68", x"d6d", x"d72", x"d76", x"d7b", x"d7f",
        x"d84", x"d88", x"d8d", x"d91", x"d96", x"d9a", x"d9f", x"da3",
        x"da8", x"dac", x"db1", x"db5", x"dba", x"dbe", x"dc2", x"dc7",
        x"dcb", x"dcf", x"dd4", x"dd8", x"ddc", x"de0", x"de5", x"de9",
        x"ded", x"df1", x"df6", x"dfa", x"dfe", x"e02", x"e06", x"e0a",
        x"e0e", x"e13", x"e17", x"e1b", x"e1f", x"e23", x"e27", x"e2b",
        x"e2f", x"e33", x"e37", x"e3b", x"e3f", x"e43", x"e46", x"e4a",
        x"e4e", x"e52", x"e56", x"e5a", x"e5e", x"e61", x"e65", x"e69",
        x"e6d", x"e70", x"e74", x"e78", x"e7b", x"e7f", x"e83", x"e86",
        x"e8a", x"e8e", x"e91", x"e95", x"e98", x"e9c", x"e9f", x"ea3",
        x"ea6", x"eaa", x"ead", x"eb1", x"eb4", x"eb8", x"ebb", x"ebf",
        x"ec2", x"ec5", x"ec9", x"ecc", x"ecf", x"ed2", x"ed6", x"ed9",
        x"edc", x"edf", x"ee3", x"ee6", x"ee9", x"eec", x"eef", x"ef2",
        x"ef6", x"ef9", x"efc", x"eff", x"f02", x"f05", x"f08", x"f0b",
        x"f0e", x"f11", x"f14", x"f17", x"f19", x"f1c", x"f1f", x"f22",
        x"f25", x"f28", x"f2a", x"f2d", x"f30", x"f33", x"f35", x"f38",
        x"f3b", x"f3e", x"f40", x"f43", x"f45", x"f48", x"f4b", x"f4d",
        x"f50", x"f52", x"f55", x"f57", x"f5a", x"f5c", x"f5f", x"f61",
        x"f64", x"f66", x"f68", x"f6b", x"f6d", x"f6f", x"f72", x"f74",
        x"f76", x"f78", x"f7b", x"f7d", x"f7f", x"f81", x"f83", x"f86",
        x"f88", x"f8a", x"f8c", x"f8e", x"f90", x"f92", x"f94", x"f96",
        x"f98", x"f9a", x"f9c", x"f9e", x"fa0", x"fa2", x"fa4", x"fa5",
        x"fa7", x"fa9", x"fab", x"fad", x"fae", x"fb0", x"fb2", x"fb3",
        x"fb5", x"fb7", x"fb8", x"fba", x"fbc", x"fbd", x"fbf", x"fc0",
        x"fc2", x"fc3", x"fc5", x"fc6", x"fc8", x"fc9", x"fcb", x"fcc",
        x"fce", x"fcf", x"fd0", x"fd2", x"fd3", x"fd4", x"fd5", x"fd7",
        x"fd8", x"fd9", x"fda", x"fdc", x"fdd", x"fde", x"fdf", x"fe0",
        x"fe1", x"fe2", x"fe3", x"fe4", x"fe5", x"fe6", x"fe7", x"fe8",
        x"fe9", x"fea", x"feb", x"fec", x"fed", x"fed", x"fee", x"fef",
        x"ff0", x"ff1", x"ff1", x"ff2", x"ff3", x"ff3", x"ff4", x"ff5",
        x"ff5", x"ff6", x"ff6", x"ff7", x"ff8", x"ff8", x"ff9", x"ff9",
        x"ffa", x"ffa", x"ffa", x"ffb", x"ffb", x"ffc", x"ffc", x"ffc",
        x"ffd", x"ffd", x"ffd", x"ffd", x"ffe", x"ffe", x"ffe", x"ffe",
        x"ffe", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ffe",
        x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffd", x"ffd", x"ffd",
        x"ffc", x"ffc", x"ffc", x"ffb", x"ffb", x"ffb", x"ffa", x"ffa",
        x"ff9", x"ff9", x"ff8", x"ff8", x"ff7", x"ff7", x"ff6", x"ff6",
        x"ff5", x"ff4", x"ff4", x"ff3", x"ff2", x"ff2", x"ff1", x"ff0",
        x"fef", x"fef", x"fee", x"fed", x"fec", x"feb", x"fea", x"fea",
        x"fe9", x"fe8", x"fe7", x"fe6", x"fe5", x"fe4", x"fe3", x"fe2",
        x"fe1", x"fdf", x"fde", x"fdd", x"fdc", x"fdb", x"fda", x"fd9",
        x"fd7", x"fd6", x"fd5", x"fd4", x"fd2", x"fd1", x"fd0", x"fce",
        x"fcd", x"fcb", x"fca", x"fc9", x"fc7", x"fc6", x"fc4", x"fc3",
        x"fc1", x"fc0", x"fbe", x"fbd", x"fbb", x"fb9", x"fb8", x"fb6",
        x"fb4", x"fb3", x"fb1", x"faf", x"fad", x"fac", x"faa", x"fa8",
        x"fa6", x"fa4", x"fa3", x"fa1", x"f9f", x"f9d", x"f9b", x"f99",
        x"f97", x"f95", x"f93", x"f91", x"f8f", x"f8d", x"f8b", x"f89",
        x"f87", x"f85", x"f82", x"f80", x"f7e", x"f7c", x"f7a", x"f77",
        x"f75", x"f73", x"f71", x"f6e", x"f6c", x"f6a", x"f67", x"f65",
        x"f62", x"f60", x"f5e", x"f5b", x"f59", x"f56", x"f54", x"f51",
        x"f4f", x"f4c", x"f49", x"f47", x"f44", x"f42", x"f3f", x"f3c",
        x"f3a", x"f37", x"f34", x"f31", x"f2f", x"f2c", x"f29", x"f26",
        x"f23", x"f21", x"f1e", x"f1b", x"f18", x"f15", x"f12", x"f0f",
        x"f0c", x"f09", x"f06", x"f03", x"f00", x"efd", x"efa", x"ef7",
        x"ef4", x"ef1", x"eee", x"eeb", x"ee7", x"ee4", x"ee1", x"ede",
        x"edb", x"ed7", x"ed4", x"ed1", x"ece", x"eca", x"ec7", x"ec4",
        x"ec0", x"ebd", x"eb9", x"eb6", x"eb3", x"eaf", x"eac", x"ea8",
        x"ea5", x"ea1", x"e9e", x"e9a", x"e97", x"e93", x"e8f", x"e8c",
        x"e88", x"e85", x"e81", x"e7d", x"e7a", x"e76", x"e72", x"e6e",
        x"e6b", x"e67", x"e63", x"e5f", x"e5c", x"e58", x"e54", x"e50",
        x"e4c", x"e48", x"e44", x"e41", x"e3d", x"e39", x"e35", x"e31",
        x"e2d", x"e29", x"e25", x"e21", x"e1d", x"e19", x"e15", x"e10",
        x"e0c", x"e08", x"e04", x"e00", x"dfc", x"df8", x"df3", x"def",
        x"deb", x"de7", x"de3", x"dde", x"dda", x"dd6", x"dd1", x"dcd",
        x"dc9", x"dc4", x"dc0", x"dbc", x"db7", x"db3", x"daf", x"daa",
        x"da6", x"da1", x"d9d", x"d98", x"d94", x"d8f", x"d8b", x"d86",
        x"d82", x"d7d", x"d78", x"d74", x"d6f", x"d6b", x"d66", x"d61",
        x"d5d", x"d58", x"d53", x"d4f", x"d4a", x"d45", x"d41", x"d3c",
        x"d37", x"d32", x"d2d", x"d29", x"d24", x"d1f", x"d1a", x"d15",
        x"d11", x"d0c", x"d07", x"d02", x"cfd", x"cf8", x"cf3", x"cee",
        x"ce9", x"ce4", x"cdf", x"cda", x"cd5", x"cd0", x"ccb", x"cc6",
        x"cc1", x"cbc", x"cb7", x"cb2", x"cad", x"ca8", x"ca3", x"c9e",
        x"c98", x"c93", x"c8e", x"c89", x"c84", x"c7f", x"c79", x"c74",
        x"c6f", x"c6a", x"c64", x"c5f", x"c5a", x"c55", x"c4f", x"c4a",
        x"c45", x"c3f", x"c3a", x"c35", x"c2f", x"c2a", x"c25", x"c1f",
        x"c1a", x"c14", x"c0f", x"c0a", x"c04", x"bff", x"bf9", x"bf4",
        x"bee", x"be9", x"be3", x"bde", x"bd8", x"bd3", x"bcd", x"bc8",
        x"bc2", x"bbd", x"bb7", x"bb2", x"bac", x"ba7", x"ba1", x"b9b",
        x"b96", x"b90", x"b8a", x"b85", x"b7f", x"b79", x"b74", x"b6e",
        x"b68", x"b63", x"b5d", x"b57", x"b52", x"b4c", x"b46", x"b40",
        x"b3b", x"b35", x"b2f", x"b29", x"b24", x"b1e", x"b18", x"b12",
        x"b0d", x"b07", x"b01", x"afb", x"af5", x"aef", x"aea", x"ae4",
        x"ade", x"ad8", x"ad2", x"acc", x"ac6", x"ac0", x"aba", x"ab5",
        x"aaf", x"aa9", x"aa3", x"a9d", x"a97", x"a91", x"a8b", x"a85",
        x"a7f", x"a79", x"a73", x"a6d", x"a67", x"a61", x"a5b", x"a55",
        x"a4f", x"a49", x"a43", x"a3d", x"a37", x"a31", x"a2b", x"a25",
        x"a1f", x"a19", x"a13", x"a0d", x"a07", x"a00", x"9fa", x"9f4",
        x"9ee", x"9e8", x"9e2", x"9dc", x"9d6", x"9d0", x"9ca", x"9c3",
        x"9bd", x"9b7", x"9b1", x"9ab", x"9a5", x"99f", x"998", x"992",
        x"98c", x"986", x"980", x"97a", x"973", x"96d", x"967", x"961",
        x"95b", x"954", x"94e", x"948", x"942", x"93c", x"935", x"92f",
        x"929", x"923", x"91d", x"916", x"910", x"90a", x"904", x"8fd",
        x"8f7", x"8f1", x"8eb", x"8e4", x"8de", x"8d8", x"8d2", x"8cb",
        x"8c5", x"8bf", x"8b9", x"8b2", x"8ac", x"8a6", x"8a0", x"899",
        x"893", x"88d", x"887", x"880", x"87a", x"874", x"86d", x"867",
        x"861", x"85b", x"854", x"84e", x"848", x"841", x"83b", x"835",
        x"82f", x"828", x"822", x"81c", x"815", x"80f", x"809", x"803",
        x"7fc", x"7f6", x"7f0", x"7ea", x"7e3", x"7dd", x"7d7", x"7d0",
        x"7ca", x"7c4", x"7be", x"7b7", x"7b1", x"7ab", x"7a4", x"79e",
        x"798", x"792", x"78b", x"785", x"77f", x"778", x"772", x"76c",
        x"766", x"75f", x"759", x"753", x"74d", x"746", x"740", x"73a",
        x"734", x"72d", x"727", x"721", x"71b", x"714", x"70e", x"708",
        x"702", x"6fb", x"6f5", x"6ef", x"6e9", x"6e2", x"6dc", x"6d6",
        x"6d0", x"6ca", x"6c3", x"6bd", x"6b7", x"6b1", x"6ab", x"6a4",
        x"69e", x"698", x"692", x"68c", x"685", x"67f", x"679", x"673",
        x"66d", x"667", x"660", x"65a", x"654", x"64e", x"648", x"642",
        x"63c", x"635", x"62f", x"629", x"623", x"61d", x"617", x"611",
        x"60b", x"605", x"5ff", x"5f8", x"5f2", x"5ec", x"5e6", x"5e0",
        x"5da", x"5d4", x"5ce", x"5c8", x"5c2", x"5bc", x"5b6", x"5b0",
        x"5aa", x"5a4", x"59e", x"598", x"592", x"58c", x"586", x"580",
        x"57a", x"574", x"56e", x"568", x"562", x"55c", x"556", x"550",
        x"54a", x"545", x"53f", x"539", x"533", x"52d", x"527", x"521",
        x"51b", x"515", x"510", x"50a", x"504", x"4fe", x"4f8", x"4f2",
        x"4ed", x"4e7", x"4e1", x"4db", x"4d6", x"4d0", x"4ca", x"4c4",
        x"4bf", x"4b9", x"4b3", x"4ad", x"4a8", x"4a2", x"49c", x"497",
        x"491", x"48b", x"486", x"480", x"47a", x"475", x"46f", x"469",
        x"464", x"45e", x"458", x"453", x"44d", x"448", x"442", x"43d",
        x"437", x"432", x"42c", x"427", x"421", x"41c", x"416", x"411",
        x"40b", x"406", x"400", x"3fb", x"3f5", x"3f0", x"3eb", x"3e5",
        x"3e0", x"3da", x"3d5", x"3d0", x"3ca", x"3c5", x"3c0", x"3ba",
        x"3b5", x"3b0", x"3aa", x"3a5", x"3a0", x"39b", x"395", x"390",
        x"38b", x"386", x"380", x"37b", x"376", x"371", x"36c", x"367",
        x"361", x"35c", x"357", x"352", x"34d", x"348", x"343", x"33e",
        x"339", x"334", x"32f", x"32a", x"325", x"320", x"31b", x"316",
        x"311", x"30c", x"307", x"302", x"2fd", x"2f8", x"2f3", x"2ee",
        x"2ea", x"2e5", x"2e0", x"2db", x"2d6", x"2d2", x"2cd", x"2c8",
        x"2c3", x"2be", x"2ba", x"2b5", x"2b0", x"2ac", x"2a7", x"2a2",
        x"29e", x"299", x"294", x"290", x"28b", x"287", x"282", x"27d",
        x"279", x"274", x"270", x"26b", x"267", x"262", x"25e", x"259",
        x"255", x"250", x"24c", x"248", x"243", x"23f", x"23b", x"236",
        x"232", x"22e", x"229", x"225", x"221", x"21c", x"218", x"214",
        x"210", x"20c", x"207", x"203", x"1ff", x"1fb", x"1f7", x"1f3",
        x"1ef", x"1ea", x"1e6", x"1e2", x"1de", x"1da", x"1d6", x"1d2",
        x"1ce", x"1ca", x"1c6", x"1c2", x"1be", x"1bb", x"1b7", x"1b3",
        x"1af", x"1ab", x"1a7", x"1a3", x"1a0", x"19c", x"198", x"194",
        x"191", x"18d", x"189", x"185", x"182", x"17e", x"17a", x"177",
        x"173", x"170", x"16c", x"168", x"165", x"161", x"15e", x"15a",
        x"157", x"153", x"150", x"14c", x"149", x"146", x"142", x"13f",
        x"13b", x"138", x"135", x"131", x"12e", x"12b", x"128", x"124",
        x"121", x"11e", x"11b", x"118", x"114", x"111", x"10e", x"10b",
        x"108", x"105", x"102", x"0ff", x"0fc", x"0f9", x"0f6", x"0f3",
        x"0f0", x"0ed", x"0ea", x"0e7", x"0e4", x"0e1", x"0de", x"0dc",
        x"0d9", x"0d6", x"0d3", x"0d0", x"0ce", x"0cb", x"0c8", x"0c5",
        x"0c3", x"0c0", x"0bd", x"0bb", x"0b8", x"0b6", x"0b3", x"0b0",
        x"0ae", x"0ab", x"0a9", x"0a6", x"0a4", x"0a1", x"09f", x"09d",
        x"09a", x"098", x"095", x"093", x"091", x"08e", x"08c", x"08a",
        x"088", x"085", x"083", x"081", x"07f", x"07d", x"07a", x"078",
        x"076", x"074", x"072", x"070", x"06e", x"06c", x"06a", x"068",
        x"066", x"064", x"062", x"060", x"05e", x"05c", x"05b", x"059",
        x"057", x"055", x"053", x"052", x"050", x"04e", x"04c", x"04b",
        x"049", x"047", x"046", x"044", x"042", x"041", x"03f", x"03e",
        x"03c", x"03b", x"039", x"038", x"036", x"035", x"034", x"032",
        x"031", x"02f", x"02e", x"02d", x"02b", x"02a", x"029", x"028",
        x"026", x"025", x"024", x"023", x"022", x"021", x"020", x"01e",
        x"01d", x"01c", x"01b", x"01a", x"019", x"018", x"017", x"016",
        x"015", x"015", x"014", x"013", x"012", x"011", x"010", x"010",
        x"00f", x"00e", x"00d", x"00d", x"00c", x"00b", x"00b", x"00a",
        x"009", x"009", x"008", x"008", x"007", x"007", x"006", x"006",
        x"005", x"005", x"004", x"004", x"004", x"003", x"003", x"003",
        x"002", x"002", x"002", x"001", x"001", x"001", x"001", x"001",
        x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
        x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"001",
        x"001", x"001", x"001", x"001", x"002", x"002", x"002", x"002",
        x"003", x"003", x"003", x"004", x"004", x"005", x"005", x"005",
        x"006", x"006", x"007", x"007", x"008", x"009", x"009", x"00a",
        x"00a", x"00b", x"00c", x"00c", x"00d", x"00e", x"00e", x"00f",
        x"010", x"011", x"012", x"012", x"013", x"014", x"015", x"016",
        x"017", x"018", x"019", x"01a", x"01b", x"01c", x"01d", x"01e",
        x"01f", x"020", x"021", x"022", x"023", x"025", x"026", x"027",
        x"028", x"02a", x"02b", x"02c", x"02d", x"02f", x"030", x"031",
        x"033", x"034", x"036", x"037", x"039", x"03a", x"03c", x"03d",
        x"03f", x"040", x"042", x"043", x"045", x"047", x"048", x"04a",
        x"04c", x"04d", x"04f", x"051", x"052", x"054", x"056", x"058",
        x"05a", x"05b", x"05d", x"05f", x"061", x"063", x"065", x"067",
        x"069", x"06b", x"06d", x"06f", x"071", x"073", x"075", x"077",
        x"079", x"07c", x"07e", x"080", x"082", x"084", x"087", x"089",
        x"08b", x"08d", x"090", x"092", x"094", x"097", x"099", x"09b",
        x"09e", x"0a0", x"0a3", x"0a5", x"0a8", x"0aa", x"0ad", x"0af",
        x"0b2", x"0b4", x"0b7", x"0ba", x"0bc", x"0bf", x"0c1", x"0c4",
        x"0c7", x"0ca", x"0cc", x"0cf", x"0d2", x"0d5", x"0d7", x"0da",
        x"0dd", x"0e0", x"0e3", x"0e6", x"0e8", x"0eb", x"0ee", x"0f1",
        x"0f4", x"0f7", x"0fa", x"0fd", x"100", x"103", x"106", x"109",
        x"10d", x"110", x"113", x"116", x"119", x"11c", x"120", x"123",
        x"126", x"129", x"12d", x"130", x"133", x"136", x"13a", x"13d",
        x"140", x"144", x"147", x"14b", x"14e", x"152", x"155", x"159",
        x"15c", x"160", x"163", x"167", x"16a", x"16e", x"171", x"175",
        x"179", x"17c", x"180", x"184", x"187", x"18b", x"18f", x"192",
        x"196", x"19a", x"19e", x"1a1", x"1a5", x"1a9", x"1ad", x"1b1",
        x"1b5", x"1b9", x"1bc", x"1c0", x"1c4", x"1c8", x"1cc", x"1d0",
        x"1d4", x"1d8", x"1dc", x"1e0", x"1e4", x"1e8", x"1ec", x"1f1",
        x"1f5", x"1f9", x"1fd", x"201", x"205", x"209", x"20e", x"212",
        x"216", x"21a", x"21f", x"223", x"227", x"22b", x"230", x"234",
        x"238", x"23d", x"241", x"245", x"24a", x"24e", x"253", x"257",
        x"25c", x"260", x"265", x"269", x"26e", x"272", x"277", x"27b",
        x"280", x"284", x"289", x"28d", x"292", x"297", x"29b", x"2a0",
        x"2a5", x"2a9", x"2ae", x"2b3", x"2b7", x"2bc", x"2c1", x"2c6",
        x"2ca", x"2cf", x"2d4", x"2d9", x"2de", x"2e2", x"2e7", x"2ec",
        x"2f1", x"2f6", x"2fb", x"300", x"304", x"309", x"30e", x"313",
        x"318", x"31d", x"322", x"327", x"32c", x"331", x"336", x"33b",
        x"340", x"345", x"34a", x"350", x"355", x"35a", x"35f", x"364",
        x"369", x"36e", x"373", x"379", x"37e", x"383", x"388", x"38d",
        x"393", x"398", x"39d", x"3a2", x"3a8", x"3ad", x"3b2", x"3b8",
        x"3bd", x"3c2", x"3c8", x"3cd", x"3d2", x"3d8", x"3dd", x"3e2",
        x"3e8", x"3ed", x"3f3", x"3f8", x"3fd", x"403", x"408", x"40e",
        x"413", x"419", x"41e", x"424", x"429", x"42f", x"434", x"43a",
        x"43f", x"445", x"44b", x"450", x"456", x"45b", x"461", x"467",
        x"46c", x"472", x"477", x"47d", x"483", x"488", x"48e", x"494",
        x"499", x"49f", x"4a5", x"4aa", x"4b0", x"4b6", x"4bc", x"4c1",
        x"4c7", x"4cd", x"4d3", x"4d8", x"4de", x"4e4", x"4ea", x"4f0",
        x"4f5", x"4fb", x"501", x"507", x"50d", x"513", x"518", x"51e",
        x"524", x"52a", x"530", x"536", x"53c", x"542", x"547", x"54d",
        x"553", x"559", x"55f", x"565", x"56b", x"571", x"577", x"57d",
        x"583", x"589", x"58f", x"595", x"59b", x"5a1", x"5a7", x"5ad",
        x"5b3", x"5b9", x"5bf", x"5c5", x"5cb", x"5d1", x"5d7", x"5dd",
        x"5e3", x"5e9", x"5ef", x"5f5", x"5fb", x"602", x"608", x"60e",
        x"614", x"61a", x"620", x"626", x"62c", x"632", x"639", x"63f",
        x"645", x"64b", x"651", x"657", x"65d", x"664", x"66a", x"670",
        x"676", x"67c", x"682", x"689", x"68f", x"695", x"69b", x"6a1",
        x"6a7", x"6ae", x"6b4", x"6ba", x"6c0", x"6c6", x"6cd", x"6d3",
        x"6d9", x"6df", x"6e6", x"6ec", x"6f2", x"6f8", x"6ff", x"705",
        x"70b", x"711", x"717", x"71e", x"724", x"72a", x"730", x"737",
        x"73d", x"743", x"749", x"750", x"756", x"75c", x"763", x"769",
        x"76f", x"775", x"77c", x"782", x"788", x"78e", x"795", x"79b",
        x"7a1", x"7a8", x"7ae", x"7b4", x"7ba", x"7c1", x"7c7", x"7cd",
        x"7d4", x"7da", x"7e0", x"7e6", x"7ed", x"7f3", x"7f9", x"800"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr,clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp,en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
