library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(11 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom;

architecture arch of rom is
    type memoria_rom is array (0 to 4095) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"002", x"004", x"006", x"008", x"00a", x"00c", x"00e", x"010",
        x"012", x"014", x"016", x"018", x"01a", x"01c", x"01e", x"020",
        x"022", x"024", x"026", x"028", x"02a", x"02c", x"02e", x"030",
        x"032", x"034", x"036", x"038", x"03a", x"03c", x"03e", x"040",
        x"042", x"044", x"046", x"048", x"04a", x"04c", x"04e", x"050",
        x"052", x"054", x"056", x"058", x"05a", x"05c", x"05e", x"060",
        x"062", x"064", x"066", x"068", x"06a", x"06c", x"06e", x"070",
        x"072", x"074", x"076", x"078", x"07a", x"07c", x"07e", x"080",
        x"082", x"084", x"086", x"088", x"08a", x"08c", x"08e", x"090",
        x"092", x"094", x"096", x"098", x"09a", x"09c", x"09e", x"0a0",
        x"0a2", x"0a4", x"0a6", x"0a8", x"0aa", x"0ac", x"0ae", x"0b0",
        x"0b2", x"0b4", x"0b6", x"0b8", x"0ba", x"0bc", x"0be", x"0c0",
        x"0c2", x"0c4", x"0c6", x"0c8", x"0ca", x"0cc", x"0ce", x"0d0",
        x"0d2", x"0d4", x"0d6", x"0d8", x"0da", x"0dc", x"0de", x"0e0",
        x"0e2", x"0e4", x"0e6", x"0e8", x"0ea", x"0ec", x"0ee", x"0f0",
        x"0f2", x"0f4", x"0f6", x"0f8", x"0fa", x"0fc", x"0fe", x"100",
        x"102", x"104", x"106", x"108", x"10a", x"10c", x"10e", x"110",
        x"112", x"114", x"116", x"118", x"11a", x"11c", x"11e", x"120",
        x"122", x"124", x"126", x"128", x"12a", x"12c", x"12e", x"130",
        x"132", x"134", x"136", x"138", x"13a", x"13c", x"13e", x"140",
        x"142", x"144", x"146", x"148", x"14a", x"14c", x"14e", x"150",
        x"152", x"154", x"156", x"158", x"15a", x"15c", x"15e", x"160",
        x"162", x"164", x"166", x"168", x"16a", x"16c", x"16e", x"170",
        x"172", x"174", x"176", x"178", x"17a", x"17c", x"17e", x"180",
        x"182", x"184", x"186", x"188", x"18a", x"18c", x"18e", x"190",
        x"192", x"194", x"196", x"198", x"19a", x"19c", x"19e", x"1a0",
        x"1a2", x"1a4", x"1a6", x"1a8", x"1aa", x"1ac", x"1ae", x"1b0",
        x"1b2", x"1b4", x"1b6", x"1b8", x"1ba", x"1bc", x"1be", x"1c0",
        x"1c2", x"1c4", x"1c6", x"1c8", x"1ca", x"1cc", x"1ce", x"1d0",
        x"1d2", x"1d4", x"1d6", x"1d8", x"1da", x"1dc", x"1de", x"1e0",
        x"1e2", x"1e4", x"1e6", x"1e8", x"1ea", x"1ec", x"1ee", x"1f0",
        x"1f2", x"1f4", x"1f6", x"1f8", x"1fa", x"1fc", x"1fe", x"200",
        x"202", x"204", x"206", x"208", x"20a", x"20c", x"20e", x"210",
        x"212", x"214", x"216", x"218", x"21a", x"21c", x"21e", x"220",
        x"222", x"224", x"226", x"228", x"22a", x"22c", x"22e", x"230",
        x"232", x"234", x"236", x"238", x"23a", x"23c", x"23e", x"240",
        x"242", x"244", x"246", x"248", x"24a", x"24c", x"24e", x"250",
        x"252", x"254", x"256", x"258", x"25a", x"25c", x"25e", x"260",
        x"262", x"264", x"266", x"268", x"26a", x"26c", x"26e", x"270",
        x"272", x"274", x"276", x"278", x"27a", x"27c", x"27e", x"280",
        x"282", x"284", x"286", x"288", x"28a", x"28c", x"28e", x"290",
        x"292", x"294", x"296", x"298", x"29a", x"29c", x"29e", x"2a0",
        x"2a2", x"2a4", x"2a6", x"2a8", x"2aa", x"2ac", x"2ae", x"2b0",
        x"2b2", x"2b4", x"2b6", x"2b8", x"2ba", x"2bc", x"2be", x"2c0",
        x"2c2", x"2c4", x"2c6", x"2c8", x"2ca", x"2cc", x"2ce", x"2d0",
        x"2d2", x"2d4", x"2d6", x"2d8", x"2da", x"2dc", x"2de", x"2e0",
        x"2e2", x"2e4", x"2e6", x"2e8", x"2ea", x"2ec", x"2ee", x"2f0",
        x"2f2", x"2f4", x"2f6", x"2f8", x"2fa", x"2fc", x"2fe", x"300",
        x"302", x"304", x"306", x"308", x"30a", x"30c", x"30e", x"310",
        x"312", x"314", x"316", x"318", x"31a", x"31c", x"31e", x"320",
        x"322", x"324", x"326", x"328", x"32a", x"32c", x"32e", x"330",
        x"332", x"334", x"336", x"338", x"33a", x"33c", x"33e", x"340",
        x"342", x"344", x"346", x"348", x"34a", x"34c", x"34e", x"350",
        x"352", x"354", x"356", x"358", x"35a", x"35c", x"35e", x"360",
        x"362", x"364", x"366", x"368", x"36a", x"36c", x"36e", x"370",
        x"372", x"374", x"376", x"378", x"37a", x"37c", x"37e", x"380",
        x"382", x"384", x"386", x"388", x"38a", x"38c", x"38e", x"390",
        x"392", x"394", x"396", x"398", x"39a", x"39c", x"39e", x"3a0",
        x"3a2", x"3a4", x"3a6", x"3a8", x"3aa", x"3ac", x"3ae", x"3b0",
        x"3b2", x"3b4", x"3b6", x"3b8", x"3ba", x"3bc", x"3be", x"3c0",
        x"3c2", x"3c4", x"3c6", x"3c8", x"3ca", x"3cc", x"3ce", x"3d0",
        x"3d2", x"3d4", x"3d6", x"3d8", x"3da", x"3dc", x"3de", x"3e0",
        x"3e2", x"3e4", x"3e6", x"3e8", x"3ea", x"3ec", x"3ee", x"3f0",
        x"3f2", x"3f4", x"3f6", x"3f8", x"3fa", x"3fc", x"3fe", x"400",
        x"402", x"404", x"406", x"408", x"40a", x"40c", x"40e", x"410",
        x"412", x"414", x"416", x"418", x"41a", x"41c", x"41e", x"420",
        x"422", x"424", x"426", x"428", x"42a", x"42c", x"42e", x"430",
        x"432", x"434", x"436", x"438", x"43a", x"43c", x"43e", x"440",
        x"442", x"444", x"446", x"448", x"44a", x"44c", x"44e", x"450",
        x"452", x"454", x"456", x"458", x"45a", x"45c", x"45e", x"460",
        x"462", x"464", x"466", x"468", x"46a", x"46c", x"46e", x"470",
        x"472", x"474", x"476", x"478", x"47a", x"47c", x"47e", x"480",
        x"482", x"484", x"486", x"488", x"48a", x"48c", x"48e", x"490",
        x"492", x"494", x"496", x"498", x"49a", x"49c", x"49e", x"4a0",
        x"4a2", x"4a4", x"4a6", x"4a8", x"4aa", x"4ac", x"4ae", x"4b0",
        x"4b2", x"4b4", x"4b6", x"4b8", x"4ba", x"4bc", x"4be", x"4c0",
        x"4c2", x"4c4", x"4c6", x"4c8", x"4ca", x"4cc", x"4ce", x"4d0",
        x"4d2", x"4d4", x"4d6", x"4d8", x"4da", x"4dc", x"4de", x"4e0",
        x"4e2", x"4e4", x"4e6", x"4e8", x"4ea", x"4ec", x"4ee", x"4f0",
        x"4f2", x"4f4", x"4f6", x"4f8", x"4fa", x"4fc", x"4fe", x"500",
        x"502", x"504", x"506", x"508", x"50a", x"50c", x"50e", x"510",
        x"512", x"514", x"516", x"518", x"51a", x"51c", x"51e", x"520",
        x"522", x"524", x"526", x"528", x"52a", x"52c", x"52e", x"530",
        x"532", x"534", x"536", x"538", x"53a", x"53c", x"53e", x"540",
        x"542", x"544", x"546", x"548", x"54a", x"54c", x"54e", x"550",
        x"552", x"554", x"556", x"558", x"55a", x"55c", x"55e", x"560",
        x"562", x"564", x"566", x"568", x"56a", x"56c", x"56e", x"570",
        x"572", x"574", x"576", x"578", x"57a", x"57c", x"57e", x"580",
        x"582", x"584", x"586", x"588", x"58a", x"58c", x"58e", x"590",
        x"592", x"594", x"596", x"598", x"59a", x"59c", x"59e", x"5a0",
        x"5a2", x"5a4", x"5a6", x"5a8", x"5aa", x"5ac", x"5ae", x"5b0",
        x"5b2", x"5b4", x"5b6", x"5b8", x"5ba", x"5bc", x"5be", x"5c0",
        x"5c2", x"5c4", x"5c6", x"5c8", x"5ca", x"5cc", x"5ce", x"5d0",
        x"5d2", x"5d4", x"5d6", x"5d8", x"5da", x"5dc", x"5de", x"5e0",
        x"5e2", x"5e4", x"5e6", x"5e8", x"5ea", x"5ec", x"5ee", x"5f0",
        x"5f2", x"5f4", x"5f6", x"5f8", x"5fa", x"5fc", x"5fe", x"600",
        x"602", x"604", x"606", x"608", x"60a", x"60c", x"60e", x"610",
        x"612", x"614", x"616", x"618", x"61a", x"61c", x"61e", x"620",
        x"622", x"624", x"626", x"628", x"62a", x"62c", x"62e", x"630",
        x"632", x"634", x"636", x"638", x"63a", x"63c", x"63e", x"640",
        x"642", x"644", x"646", x"648", x"64a", x"64c", x"64e", x"650",
        x"652", x"654", x"656", x"658", x"65a", x"65c", x"65e", x"660",
        x"662", x"664", x"666", x"668", x"66a", x"66c", x"66e", x"670",
        x"672", x"674", x"676", x"678", x"67a", x"67c", x"67e", x"680",
        x"682", x"684", x"686", x"688", x"68a", x"68c", x"68e", x"690",
        x"692", x"694", x"696", x"698", x"69a", x"69c", x"69e", x"6a0",
        x"6a2", x"6a4", x"6a6", x"6a8", x"6aa", x"6ac", x"6ae", x"6b0",
        x"6b2", x"6b4", x"6b6", x"6b8", x"6ba", x"6bc", x"6be", x"6c0",
        x"6c2", x"6c4", x"6c6", x"6c8", x"6ca", x"6cc", x"6ce", x"6d0",
        x"6d2", x"6d4", x"6d6", x"6d8", x"6da", x"6dc", x"6de", x"6e0",
        x"6e2", x"6e4", x"6e6", x"6e8", x"6ea", x"6ec", x"6ee", x"6f0",
        x"6f2", x"6f4", x"6f6", x"6f8", x"6fa", x"6fc", x"6fe", x"700",
        x"702", x"704", x"706", x"708", x"70a", x"70c", x"70e", x"710",
        x"712", x"714", x"716", x"718", x"71a", x"71c", x"71e", x"720",
        x"722", x"724", x"726", x"728", x"72a", x"72c", x"72e", x"730",
        x"732", x"734", x"736", x"738", x"73a", x"73c", x"73e", x"740",
        x"742", x"744", x"746", x"748", x"74a", x"74c", x"74e", x"750",
        x"752", x"754", x"756", x"758", x"75a", x"75c", x"75e", x"760",
        x"762", x"764", x"766", x"768", x"76a", x"76c", x"76e", x"770",
        x"772", x"774", x"776", x"778", x"77a", x"77c", x"77e", x"780",
        x"782", x"784", x"786", x"788", x"78a", x"78c", x"78e", x"790",
        x"792", x"794", x"796", x"798", x"79a", x"79c", x"79e", x"7a0",
        x"7a2", x"7a4", x"7a6", x"7a8", x"7aa", x"7ac", x"7ae", x"7b0",
        x"7b2", x"7b4", x"7b6", x"7b8", x"7ba", x"7bc", x"7be", x"7c0",
        x"7c2", x"7c4", x"7c6", x"7c8", x"7ca", x"7cc", x"7ce", x"7d0",
        x"7d2", x"7d4", x"7d6", x"7d8", x"7da", x"7dc", x"7de", x"7e0",
        x"7e2", x"7e4", x"7e6", x"7e8", x"7ea", x"7ec", x"7ee", x"7f0",
        x"7f2", x"7f4", x"7f6", x"7f8", x"7fa", x"7fc", x"7fe", x"800",
        x"801", x"803", x"805", x"807", x"809", x"80b", x"80d", x"80f",
        x"811", x"813", x"815", x"817", x"819", x"81b", x"81d", x"81f",
        x"821", x"823", x"825", x"827", x"829", x"82b", x"82d", x"82f",
        x"831", x"833", x"835", x"837", x"839", x"83b", x"83d", x"83f",
        x"841", x"843", x"845", x"847", x"849", x"84b", x"84d", x"84f",
        x"851", x"853", x"855", x"857", x"859", x"85b", x"85d", x"85f",
        x"861", x"863", x"865", x"867", x"869", x"86b", x"86d", x"86f",
        x"871", x"873", x"875", x"877", x"879", x"87b", x"87d", x"87f",
        x"881", x"883", x"885", x"887", x"889", x"88b", x"88d", x"88f",
        x"891", x"893", x"895", x"897", x"899", x"89b", x"89d", x"89f",
        x"8a1", x"8a3", x"8a5", x"8a7", x"8a9", x"8ab", x"8ad", x"8af",
        x"8b1", x"8b3", x"8b5", x"8b7", x"8b9", x"8bb", x"8bd", x"8bf",
        x"8c1", x"8c3", x"8c5", x"8c7", x"8c9", x"8cb", x"8cd", x"8cf",
        x"8d1", x"8d3", x"8d5", x"8d7", x"8d9", x"8db", x"8dd", x"8df",
        x"8e1", x"8e3", x"8e5", x"8e7", x"8e9", x"8eb", x"8ed", x"8ef",
        x"8f1", x"8f3", x"8f5", x"8f7", x"8f9", x"8fb", x"8fd", x"8ff",
        x"901", x"903", x"905", x"907", x"909", x"90b", x"90d", x"90f",
        x"911", x"913", x"915", x"917", x"919", x"91b", x"91d", x"91f",
        x"921", x"923", x"925", x"927", x"929", x"92b", x"92d", x"92f",
        x"931", x"933", x"935", x"937", x"939", x"93b", x"93d", x"93f",
        x"941", x"943", x"945", x"947", x"949", x"94b", x"94d", x"94f",
        x"951", x"953", x"955", x"957", x"959", x"95b", x"95d", x"95f",
        x"961", x"963", x"965", x"967", x"969", x"96b", x"96d", x"96f",
        x"971", x"973", x"975", x"977", x"979", x"97b", x"97d", x"97f",
        x"981", x"983", x"985", x"987", x"989", x"98b", x"98d", x"98f",
        x"991", x"993", x"995", x"997", x"999", x"99b", x"99d", x"99f",
        x"9a1", x"9a3", x"9a5", x"9a7", x"9a9", x"9ab", x"9ad", x"9af",
        x"9b1", x"9b3", x"9b5", x"9b7", x"9b9", x"9bb", x"9bd", x"9bf",
        x"9c1", x"9c3", x"9c5", x"9c7", x"9c9", x"9cb", x"9cd", x"9cf",
        x"9d1", x"9d3", x"9d5", x"9d7", x"9d9", x"9db", x"9dd", x"9df",
        x"9e1", x"9e3", x"9e5", x"9e7", x"9e9", x"9eb", x"9ed", x"9ef",
        x"9f1", x"9f3", x"9f5", x"9f7", x"9f9", x"9fb", x"9fd", x"9ff",
        x"a01", x"a03", x"a05", x"a07", x"a09", x"a0b", x"a0d", x"a0f",
        x"a11", x"a13", x"a15", x"a17", x"a19", x"a1b", x"a1d", x"a1f",
        x"a21", x"a23", x"a25", x"a27", x"a29", x"a2b", x"a2d", x"a2f",
        x"a31", x"a33", x"a35", x"a37", x"a39", x"a3b", x"a3d", x"a3f",
        x"a41", x"a43", x"a45", x"a47", x"a49", x"a4b", x"a4d", x"a4f",
        x"a51", x"a53", x"a55", x"a57", x"a59", x"a5b", x"a5d", x"a5f",
        x"a61", x"a63", x"a65", x"a67", x"a69", x"a6b", x"a6d", x"a6f",
        x"a71", x"a73", x"a75", x"a77", x"a79", x"a7b", x"a7d", x"a7f",
        x"a81", x"a83", x"a85", x"a87", x"a89", x"a8b", x"a8d", x"a8f",
        x"a91", x"a93", x"a95", x"a97", x"a99", x"a9b", x"a9d", x"a9f",
        x"aa1", x"aa3", x"aa5", x"aa7", x"aa9", x"aab", x"aad", x"aaf",
        x"ab1", x"ab3", x"ab5", x"ab7", x"ab9", x"abb", x"abd", x"abf",
        x"ac1", x"ac3", x"ac5", x"ac7", x"ac9", x"acb", x"acd", x"acf",
        x"ad1", x"ad3", x"ad5", x"ad7", x"ad9", x"adb", x"add", x"adf",
        x"ae1", x"ae3", x"ae5", x"ae7", x"ae9", x"aeb", x"aed", x"aef",
        x"af1", x"af3", x"af5", x"af7", x"af9", x"afb", x"afd", x"aff",
        x"b01", x"b03", x"b05", x"b07", x"b09", x"b0b", x"b0d", x"b0f",
        x"b11", x"b13", x"b15", x"b17", x"b19", x"b1b", x"b1d", x"b1f",
        x"b21", x"b23", x"b25", x"b27", x"b29", x"b2b", x"b2d", x"b2f",
        x"b31", x"b33", x"b35", x"b37", x"b39", x"b3b", x"b3d", x"b3f",
        x"b41", x"b43", x"b45", x"b47", x"b49", x"b4b", x"b4d", x"b4f",
        x"b51", x"b53", x"b55", x"b57", x"b59", x"b5b", x"b5d", x"b5f",
        x"b61", x"b63", x"b65", x"b67", x"b69", x"b6b", x"b6d", x"b6f",
        x"b71", x"b73", x"b75", x"b77", x"b79", x"b7b", x"b7d", x"b7f",
        x"b81", x"b83", x"b85", x"b87", x"b89", x"b8b", x"b8d", x"b8f",
        x"b91", x"b93", x"b95", x"b97", x"b99", x"b9b", x"b9d", x"b9f",
        x"ba1", x"ba3", x"ba5", x"ba7", x"ba9", x"bab", x"bad", x"baf",
        x"bb1", x"bb3", x"bb5", x"bb7", x"bb9", x"bbb", x"bbd", x"bbf",
        x"bc1", x"bc3", x"bc5", x"bc7", x"bc9", x"bcb", x"bcd", x"bcf",
        x"bd1", x"bd3", x"bd5", x"bd7", x"bd9", x"bdb", x"bdd", x"bdf",
        x"be1", x"be3", x"be5", x"be7", x"be9", x"beb", x"bed", x"bef",
        x"bf1", x"bf3", x"bf5", x"bf7", x"bf9", x"bfb", x"bfd", x"bff",
        x"c01", x"c03", x"c05", x"c07", x"c09", x"c0b", x"c0d", x"c0f",
        x"c11", x"c13", x"c15", x"c17", x"c19", x"c1b", x"c1d", x"c1f",
        x"c21", x"c23", x"c25", x"c27", x"c29", x"c2b", x"c2d", x"c2f",
        x"c31", x"c33", x"c35", x"c37", x"c39", x"c3b", x"c3d", x"c3f",
        x"c41", x"c43", x"c45", x"c47", x"c49", x"c4b", x"c4d", x"c4f",
        x"c51", x"c53", x"c55", x"c57", x"c59", x"c5b", x"c5d", x"c5f",
        x"c61", x"c63", x"c65", x"c67", x"c69", x"c6b", x"c6d", x"c6f",
        x"c71", x"c73", x"c75", x"c77", x"c79", x"c7b", x"c7d", x"c7f",
        x"c81", x"c83", x"c85", x"c87", x"c89", x"c8b", x"c8d", x"c8f",
        x"c91", x"c93", x"c95", x"c97", x"c99", x"c9b", x"c9d", x"c9f",
        x"ca1", x"ca3", x"ca5", x"ca7", x"ca9", x"cab", x"cad", x"caf",
        x"cb1", x"cb3", x"cb5", x"cb7", x"cb9", x"cbb", x"cbd", x"cbf",
        x"cc1", x"cc3", x"cc5", x"cc7", x"cc9", x"ccb", x"ccd", x"ccf",
        x"cd1", x"cd3", x"cd5", x"cd7", x"cd9", x"cdb", x"cdd", x"cdf",
        x"ce1", x"ce3", x"ce5", x"ce7", x"ce9", x"ceb", x"ced", x"cef",
        x"cf1", x"cf3", x"cf5", x"cf7", x"cf9", x"cfb", x"cfd", x"cff",
        x"d01", x"d03", x"d05", x"d07", x"d09", x"d0b", x"d0d", x"d0f",
        x"d11", x"d13", x"d15", x"d17", x"d19", x"d1b", x"d1d", x"d1f",
        x"d21", x"d23", x"d25", x"d27", x"d29", x"d2b", x"d2d", x"d2f",
        x"d31", x"d33", x"d35", x"d37", x"d39", x"d3b", x"d3d", x"d3f",
        x"d41", x"d43", x"d45", x"d47", x"d49", x"d4b", x"d4d", x"d4f",
        x"d51", x"d53", x"d55", x"d57", x"d59", x"d5b", x"d5d", x"d5f",
        x"d61", x"d63", x"d65", x"d67", x"d69", x"d6b", x"d6d", x"d6f",
        x"d71", x"d73", x"d75", x"d77", x"d79", x"d7b", x"d7d", x"d7f",
        x"d81", x"d83", x"d85", x"d87", x"d89", x"d8b", x"d8d", x"d8f",
        x"d91", x"d93", x"d95", x"d97", x"d99", x"d9b", x"d9d", x"d9f",
        x"da1", x"da3", x"da5", x"da7", x"da9", x"dab", x"dad", x"daf",
        x"db1", x"db3", x"db5", x"db7", x"db9", x"dbb", x"dbd", x"dbf",
        x"dc1", x"dc3", x"dc5", x"dc7", x"dc9", x"dcb", x"dcd", x"dcf",
        x"dd1", x"dd3", x"dd5", x"dd7", x"dd9", x"ddb", x"ddd", x"ddf",
        x"de1", x"de3", x"de5", x"de7", x"de9", x"deb", x"ded", x"def",
        x"df1", x"df3", x"df5", x"df7", x"df9", x"dfb", x"dfd", x"dff",
        x"e01", x"e03", x"e05", x"e07", x"e09", x"e0b", x"e0d", x"e0f",
        x"e11", x"e13", x"e15", x"e17", x"e19", x"e1b", x"e1d", x"e1f",
        x"e21", x"e23", x"e25", x"e27", x"e29", x"e2b", x"e2d", x"e2f",
        x"e31", x"e33", x"e35", x"e37", x"e39", x"e3b", x"e3d", x"e3f",
        x"e41", x"e43", x"e45", x"e47", x"e49", x"e4b", x"e4d", x"e4f",
        x"e51", x"e53", x"e55", x"e57", x"e59", x"e5b", x"e5d", x"e5f",
        x"e61", x"e63", x"e65", x"e67", x"e69", x"e6b", x"e6d", x"e6f",
        x"e71", x"e73", x"e75", x"e77", x"e79", x"e7b", x"e7d", x"e7f",
        x"e81", x"e83", x"e85", x"e87", x"e89", x"e8b", x"e8d", x"e8f",
        x"e91", x"e93", x"e95", x"e97", x"e99", x"e9b", x"e9d", x"e9f",
        x"ea1", x"ea3", x"ea5", x"ea7", x"ea9", x"eab", x"ead", x"eaf",
        x"eb1", x"eb3", x"eb5", x"eb7", x"eb9", x"ebb", x"ebd", x"ebf",
        x"ec1", x"ec3", x"ec5", x"ec7", x"ec9", x"ecb", x"ecd", x"ecf",
        x"ed1", x"ed3", x"ed5", x"ed7", x"ed9", x"edb", x"edd", x"edf",
        x"ee1", x"ee3", x"ee5", x"ee7", x"ee9", x"eeb", x"eed", x"eef",
        x"ef1", x"ef3", x"ef5", x"ef7", x"ef9", x"efb", x"efd", x"eff",
        x"f01", x"f03", x"f05", x"f07", x"f09", x"f0b", x"f0d", x"f0f",
        x"f11", x"f13", x"f15", x"f17", x"f19", x"f1b", x"f1d", x"f1f",
        x"f21", x"f23", x"f25", x"f27", x"f29", x"f2b", x"f2d", x"f2f",
        x"f31", x"f33", x"f35", x"f37", x"f39", x"f3b", x"f3d", x"f3f",
        x"f41", x"f43", x"f45", x"f47", x"f49", x"f4b", x"f4d", x"f4f",
        x"f51", x"f53", x"f55", x"f57", x"f59", x"f5b", x"f5d", x"f5f",
        x"f61", x"f63", x"f65", x"f67", x"f69", x"f6b", x"f6d", x"f6f",
        x"f71", x"f73", x"f75", x"f77", x"f79", x"f7b", x"f7d", x"f7f",
        x"f81", x"f83", x"f85", x"f87", x"f89", x"f8b", x"f8d", x"f8f",
        x"f91", x"f93", x"f95", x"f97", x"f99", x"f9b", x"f9d", x"f9f",
        x"fa1", x"fa3", x"fa5", x"fa7", x"fa9", x"fab", x"fad", x"faf",
        x"fb1", x"fb3", x"fb5", x"fb7", x"fb9", x"fbb", x"fbd", x"fbf",
        x"fc1", x"fc3", x"fc5", x"fc7", x"fc9", x"fcb", x"fcd", x"fcf",
        x"fd1", x"fd3", x"fd5", x"fd7", x"fd9", x"fdb", x"fdd", x"fdf",
        x"fe1", x"fe3", x"fe5", x"fe7", x"fe9", x"feb", x"fed", x"fef",
        x"ff1", x"ff3", x"ff5", x"ff7", x"ff9", x"ffb", x"ffd", x"fff",
        x"ffd", x"ffb", x"ff9", x"ff7", x"ff5", x"ff3", x"ff1", x"fef",
        x"fed", x"feb", x"fe9", x"fe7", x"fe5", x"fe3", x"fe1", x"fdf",
        x"fdd", x"fdb", x"fd9", x"fd7", x"fd5", x"fd3", x"fd1", x"fcf",
        x"fcd", x"fcb", x"fc9", x"fc7", x"fc5", x"fc3", x"fc1", x"fbf",
        x"fbd", x"fbb", x"fb9", x"fb7", x"fb5", x"fb3", x"fb1", x"faf",
        x"fad", x"fab", x"fa9", x"fa7", x"fa5", x"fa3", x"fa1", x"f9f",
        x"f9d", x"f9b", x"f99", x"f97", x"f95", x"f93", x"f91", x"f8f",
        x"f8d", x"f8b", x"f89", x"f87", x"f85", x"f83", x"f81", x"f7f",
        x"f7d", x"f7b", x"f79", x"f77", x"f75", x"f73", x"f71", x"f6f",
        x"f6d", x"f6b", x"f69", x"f67", x"f65", x"f63", x"f61", x"f5f",
        x"f5d", x"f5b", x"f59", x"f57", x"f55", x"f53", x"f51", x"f4f",
        x"f4d", x"f4b", x"f49", x"f47", x"f45", x"f43", x"f41", x"f3f",
        x"f3d", x"f3b", x"f39", x"f37", x"f35", x"f33", x"f31", x"f2f",
        x"f2d", x"f2b", x"f29", x"f27", x"f25", x"f23", x"f21", x"f1f",
        x"f1d", x"f1b", x"f19", x"f17", x"f15", x"f13", x"f11", x"f0f",
        x"f0d", x"f0b", x"f09", x"f07", x"f05", x"f03", x"f01", x"eff",
        x"efd", x"efb", x"ef9", x"ef7", x"ef5", x"ef3", x"ef1", x"eef",
        x"eed", x"eeb", x"ee9", x"ee7", x"ee5", x"ee3", x"ee1", x"edf",
        x"edd", x"edb", x"ed9", x"ed7", x"ed5", x"ed3", x"ed1", x"ecf",
        x"ecd", x"ecb", x"ec9", x"ec7", x"ec5", x"ec3", x"ec1", x"ebf",
        x"ebd", x"ebb", x"eb9", x"eb7", x"eb5", x"eb3", x"eb1", x"eaf",
        x"ead", x"eab", x"ea9", x"ea7", x"ea5", x"ea3", x"ea1", x"e9f",
        x"e9d", x"e9b", x"e99", x"e97", x"e95", x"e93", x"e91", x"e8f",
        x"e8d", x"e8b", x"e89", x"e87", x"e85", x"e83", x"e81", x"e7f",
        x"e7d", x"e7b", x"e79", x"e77", x"e75", x"e73", x"e71", x"e6f",
        x"e6d", x"e6b", x"e69", x"e67", x"e65", x"e63", x"e61", x"e5f",
        x"e5d", x"e5b", x"e59", x"e57", x"e55", x"e53", x"e51", x"e4f",
        x"e4d", x"e4b", x"e49", x"e47", x"e45", x"e43", x"e41", x"e3f",
        x"e3d", x"e3b", x"e39", x"e37", x"e35", x"e33", x"e31", x"e2f",
        x"e2d", x"e2b", x"e29", x"e27", x"e25", x"e23", x"e21", x"e1f",
        x"e1d", x"e1b", x"e19", x"e17", x"e15", x"e13", x"e11", x"e0f",
        x"e0d", x"e0b", x"e09", x"e07", x"e05", x"e03", x"e01", x"dff",
        x"dfd", x"dfb", x"df9", x"df7", x"df5", x"df3", x"df1", x"def",
        x"ded", x"deb", x"de9", x"de7", x"de5", x"de3", x"de1", x"ddf",
        x"ddd", x"ddb", x"dd9", x"dd7", x"dd5", x"dd3", x"dd1", x"dcf",
        x"dcd", x"dcb", x"dc9", x"dc7", x"dc5", x"dc3", x"dc1", x"dbf",
        x"dbd", x"dbb", x"db9", x"db7", x"db5", x"db3", x"db1", x"daf",
        x"dad", x"dab", x"da9", x"da7", x"da5", x"da3", x"da1", x"d9f",
        x"d9d", x"d9b", x"d99", x"d97", x"d95", x"d93", x"d91", x"d8f",
        x"d8d", x"d8b", x"d89", x"d87", x"d85", x"d83", x"d81", x"d7f",
        x"d7d", x"d7b", x"d79", x"d77", x"d75", x"d73", x"d71", x"d6f",
        x"d6d", x"d6b", x"d69", x"d67", x"d65", x"d63", x"d61", x"d5f",
        x"d5d", x"d5b", x"d59", x"d57", x"d55", x"d53", x"d51", x"d4f",
        x"d4d", x"d4b", x"d49", x"d47", x"d45", x"d43", x"d41", x"d3f",
        x"d3d", x"d3b", x"d39", x"d37", x"d35", x"d33", x"d31", x"d2f",
        x"d2d", x"d2b", x"d29", x"d27", x"d25", x"d23", x"d21", x"d1f",
        x"d1d", x"d1b", x"d19", x"d17", x"d15", x"d13", x"d11", x"d0f",
        x"d0d", x"d0b", x"d09", x"d07", x"d05", x"d03", x"d01", x"cff",
        x"cfd", x"cfb", x"cf9", x"cf7", x"cf5", x"cf3", x"cf1", x"cef",
        x"ced", x"ceb", x"ce9", x"ce7", x"ce5", x"ce3", x"ce1", x"cdf",
        x"cdd", x"cdb", x"cd9", x"cd7", x"cd5", x"cd3", x"cd1", x"ccf",
        x"ccd", x"ccb", x"cc9", x"cc7", x"cc5", x"cc3", x"cc1", x"cbf",
        x"cbd", x"cbb", x"cb9", x"cb7", x"cb5", x"cb3", x"cb1", x"caf",
        x"cad", x"cab", x"ca9", x"ca7", x"ca5", x"ca3", x"ca1", x"c9f",
        x"c9d", x"c9b", x"c99", x"c97", x"c95", x"c93", x"c91", x"c8f",
        x"c8d", x"c8b", x"c89", x"c87", x"c85", x"c83", x"c81", x"c7f",
        x"c7d", x"c7b", x"c79", x"c77", x"c75", x"c73", x"c71", x"c6f",
        x"c6d", x"c6b", x"c69", x"c67", x"c65", x"c63", x"c61", x"c5f",
        x"c5d", x"c5b", x"c59", x"c57", x"c55", x"c53", x"c51", x"c4f",
        x"c4d", x"c4b", x"c49", x"c47", x"c45", x"c43", x"c41", x"c3f",
        x"c3d", x"c3b", x"c39", x"c37", x"c35", x"c33", x"c31", x"c2f",
        x"c2d", x"c2b", x"c29", x"c27", x"c25", x"c23", x"c21", x"c1f",
        x"c1d", x"c1b", x"c19", x"c17", x"c15", x"c13", x"c11", x"c0f",
        x"c0d", x"c0b", x"c09", x"c07", x"c05", x"c03", x"c01", x"bff",
        x"bfd", x"bfb", x"bf9", x"bf7", x"bf5", x"bf3", x"bf1", x"bef",
        x"bed", x"beb", x"be9", x"be7", x"be5", x"be3", x"be1", x"bdf",
        x"bdd", x"bdb", x"bd9", x"bd7", x"bd5", x"bd3", x"bd1", x"bcf",
        x"bcd", x"bcb", x"bc9", x"bc7", x"bc5", x"bc3", x"bc1", x"bbf",
        x"bbd", x"bbb", x"bb9", x"bb7", x"bb5", x"bb3", x"bb1", x"baf",
        x"bad", x"bab", x"ba9", x"ba7", x"ba5", x"ba3", x"ba1", x"b9f",
        x"b9d", x"b9b", x"b99", x"b97", x"b95", x"b93", x"b91", x"b8f",
        x"b8d", x"b8b", x"b89", x"b87", x"b85", x"b83", x"b81", x"b7f",
        x"b7d", x"b7b", x"b79", x"b77", x"b75", x"b73", x"b71", x"b6f",
        x"b6d", x"b6b", x"b69", x"b67", x"b65", x"b63", x"b61", x"b5f",
        x"b5d", x"b5b", x"b59", x"b57", x"b55", x"b53", x"b51", x"b4f",
        x"b4d", x"b4b", x"b49", x"b47", x"b45", x"b43", x"b41", x"b3f",
        x"b3d", x"b3b", x"b39", x"b37", x"b35", x"b33", x"b31", x"b2f",
        x"b2d", x"b2b", x"b29", x"b27", x"b25", x"b23", x"b21", x"b1f",
        x"b1d", x"b1b", x"b19", x"b17", x"b15", x"b13", x"b11", x"b0f",
        x"b0d", x"b0b", x"b09", x"b07", x"b05", x"b03", x"b01", x"aff",
        x"afd", x"afb", x"af9", x"af7", x"af5", x"af3", x"af1", x"aef",
        x"aed", x"aeb", x"ae9", x"ae7", x"ae5", x"ae3", x"ae1", x"adf",
        x"add", x"adb", x"ad9", x"ad7", x"ad5", x"ad3", x"ad1", x"acf",
        x"acd", x"acb", x"ac9", x"ac7", x"ac5", x"ac3", x"ac1", x"abf",
        x"abd", x"abb", x"ab9", x"ab7", x"ab5", x"ab3", x"ab1", x"aaf",
        x"aad", x"aab", x"aa9", x"aa7", x"aa5", x"aa3", x"aa1", x"a9f",
        x"a9d", x"a9b", x"a99", x"a97", x"a95", x"a93", x"a91", x"a8f",
        x"a8d", x"a8b", x"a89", x"a87", x"a85", x"a83", x"a81", x"a7f",
        x"a7d", x"a7b", x"a79", x"a77", x"a75", x"a73", x"a71", x"a6f",
        x"a6d", x"a6b", x"a69", x"a67", x"a65", x"a63", x"a61", x"a5f",
        x"a5d", x"a5b", x"a59", x"a57", x"a55", x"a53", x"a51", x"a4f",
        x"a4d", x"a4b", x"a49", x"a47", x"a45", x"a43", x"a41", x"a3f",
        x"a3d", x"a3b", x"a39", x"a37", x"a35", x"a33", x"a31", x"a2f",
        x"a2d", x"a2b", x"a29", x"a27", x"a25", x"a23", x"a21", x"a1f",
        x"a1d", x"a1b", x"a19", x"a17", x"a15", x"a13", x"a11", x"a0f",
        x"a0d", x"a0b", x"a09", x"a07", x"a05", x"a03", x"a01", x"9ff",
        x"9fd", x"9fb", x"9f9", x"9f7", x"9f5", x"9f3", x"9f1", x"9ef",
        x"9ed", x"9eb", x"9e9", x"9e7", x"9e5", x"9e3", x"9e1", x"9df",
        x"9dd", x"9db", x"9d9", x"9d7", x"9d5", x"9d3", x"9d1", x"9cf",
        x"9cd", x"9cb", x"9c9", x"9c7", x"9c5", x"9c3", x"9c1", x"9bf",
        x"9bd", x"9bb", x"9b9", x"9b7", x"9b5", x"9b3", x"9b1", x"9af",
        x"9ad", x"9ab", x"9a9", x"9a7", x"9a5", x"9a3", x"9a1", x"99f",
        x"99d", x"99b", x"999", x"997", x"995", x"993", x"991", x"98f",
        x"98d", x"98b", x"989", x"987", x"985", x"983", x"981", x"97f",
        x"97d", x"97b", x"979", x"977", x"975", x"973", x"971", x"96f",
        x"96d", x"96b", x"969", x"967", x"965", x"963", x"961", x"95f",
        x"95d", x"95b", x"959", x"957", x"955", x"953", x"951", x"94f",
        x"94d", x"94b", x"949", x"947", x"945", x"943", x"941", x"93f",
        x"93d", x"93b", x"939", x"937", x"935", x"933", x"931", x"92f",
        x"92d", x"92b", x"929", x"927", x"925", x"923", x"921", x"91f",
        x"91d", x"91b", x"919", x"917", x"915", x"913", x"911", x"90f",
        x"90d", x"90b", x"909", x"907", x"905", x"903", x"901", x"8ff",
        x"8fd", x"8fb", x"8f9", x"8f7", x"8f5", x"8f3", x"8f1", x"8ef",
        x"8ed", x"8eb", x"8e9", x"8e7", x"8e5", x"8e3", x"8e1", x"8df",
        x"8dd", x"8db", x"8d9", x"8d7", x"8d5", x"8d3", x"8d1", x"8cf",
        x"8cd", x"8cb", x"8c9", x"8c7", x"8c5", x"8c3", x"8c1", x"8bf",
        x"8bd", x"8bb", x"8b9", x"8b7", x"8b5", x"8b3", x"8b1", x"8af",
        x"8ad", x"8ab", x"8a9", x"8a7", x"8a5", x"8a3", x"8a1", x"89f",
        x"89d", x"89b", x"899", x"897", x"895", x"893", x"891", x"88f",
        x"88d", x"88b", x"889", x"887", x"885", x"883", x"881", x"87f",
        x"87d", x"87b", x"879", x"877", x"875", x"873", x"871", x"86f",
        x"86d", x"86b", x"869", x"867", x"865", x"863", x"861", x"85f",
        x"85d", x"85b", x"859", x"857", x"855", x"853", x"851", x"84f",
        x"84d", x"84b", x"849", x"847", x"845", x"843", x"841", x"83f",
        x"83d", x"83b", x"839", x"837", x"835", x"833", x"831", x"82f",
        x"82d", x"82b", x"829", x"827", x"825", x"823", x"821", x"81f",
        x"81d", x"81b", x"819", x"817", x"815", x"813", x"811", x"80f",
        x"80d", x"80b", x"809", x"807", x"805", x"803", x"801", x"800",
        x"7fe", x"7fc", x"7fa", x"7f8", x"7f6", x"7f4", x"7f2", x"7f0",
        x"7ee", x"7ec", x"7ea", x"7e8", x"7e6", x"7e4", x"7e2", x"7e0",
        x"7de", x"7dc", x"7da", x"7d8", x"7d6", x"7d4", x"7d2", x"7d0",
        x"7ce", x"7cc", x"7ca", x"7c8", x"7c6", x"7c4", x"7c2", x"7c0",
        x"7be", x"7bc", x"7ba", x"7b8", x"7b6", x"7b4", x"7b2", x"7b0",
        x"7ae", x"7ac", x"7aa", x"7a8", x"7a6", x"7a4", x"7a2", x"7a0",
        x"79e", x"79c", x"79a", x"798", x"796", x"794", x"792", x"790",
        x"78e", x"78c", x"78a", x"788", x"786", x"784", x"782", x"780",
        x"77e", x"77c", x"77a", x"778", x"776", x"774", x"772", x"770",
        x"76e", x"76c", x"76a", x"768", x"766", x"764", x"762", x"760",
        x"75e", x"75c", x"75a", x"758", x"756", x"754", x"752", x"750",
        x"74e", x"74c", x"74a", x"748", x"746", x"744", x"742", x"740",
        x"73e", x"73c", x"73a", x"738", x"736", x"734", x"732", x"730",
        x"72e", x"72c", x"72a", x"728", x"726", x"724", x"722", x"720",
        x"71e", x"71c", x"71a", x"718", x"716", x"714", x"712", x"710",
        x"70e", x"70c", x"70a", x"708", x"706", x"704", x"702", x"700",
        x"6fe", x"6fc", x"6fa", x"6f8", x"6f6", x"6f4", x"6f2", x"6f0",
        x"6ee", x"6ec", x"6ea", x"6e8", x"6e6", x"6e4", x"6e2", x"6e0",
        x"6de", x"6dc", x"6da", x"6d8", x"6d6", x"6d4", x"6d2", x"6d0",
        x"6ce", x"6cc", x"6ca", x"6c8", x"6c6", x"6c4", x"6c2", x"6c0",
        x"6be", x"6bc", x"6ba", x"6b8", x"6b6", x"6b4", x"6b2", x"6b0",
        x"6ae", x"6ac", x"6aa", x"6a8", x"6a6", x"6a4", x"6a2", x"6a0",
        x"69e", x"69c", x"69a", x"698", x"696", x"694", x"692", x"690",
        x"68e", x"68c", x"68a", x"688", x"686", x"684", x"682", x"680",
        x"67e", x"67c", x"67a", x"678", x"676", x"674", x"672", x"670",
        x"66e", x"66c", x"66a", x"668", x"666", x"664", x"662", x"660",
        x"65e", x"65c", x"65a", x"658", x"656", x"654", x"652", x"650",
        x"64e", x"64c", x"64a", x"648", x"646", x"644", x"642", x"640",
        x"63e", x"63c", x"63a", x"638", x"636", x"634", x"632", x"630",
        x"62e", x"62c", x"62a", x"628", x"626", x"624", x"622", x"620",
        x"61e", x"61c", x"61a", x"618", x"616", x"614", x"612", x"610",
        x"60e", x"60c", x"60a", x"608", x"606", x"604", x"602", x"600",
        x"5fe", x"5fc", x"5fa", x"5f8", x"5f6", x"5f4", x"5f2", x"5f0",
        x"5ee", x"5ec", x"5ea", x"5e8", x"5e6", x"5e4", x"5e2", x"5e0",
        x"5de", x"5dc", x"5da", x"5d8", x"5d6", x"5d4", x"5d2", x"5d0",
        x"5ce", x"5cc", x"5ca", x"5c8", x"5c6", x"5c4", x"5c2", x"5c0",
        x"5be", x"5bc", x"5ba", x"5b8", x"5b6", x"5b4", x"5b2", x"5b0",
        x"5ae", x"5ac", x"5aa", x"5a8", x"5a6", x"5a4", x"5a2", x"5a0",
        x"59e", x"59c", x"59a", x"598", x"596", x"594", x"592", x"590",
        x"58e", x"58c", x"58a", x"588", x"586", x"584", x"582", x"580",
        x"57e", x"57c", x"57a", x"578", x"576", x"574", x"572", x"570",
        x"56e", x"56c", x"56a", x"568", x"566", x"564", x"562", x"560",
        x"55e", x"55c", x"55a", x"558", x"556", x"554", x"552", x"550",
        x"54e", x"54c", x"54a", x"548", x"546", x"544", x"542", x"540",
        x"53e", x"53c", x"53a", x"538", x"536", x"534", x"532", x"530",
        x"52e", x"52c", x"52a", x"528", x"526", x"524", x"522", x"520",
        x"51e", x"51c", x"51a", x"518", x"516", x"514", x"512", x"510",
        x"50e", x"50c", x"50a", x"508", x"506", x"504", x"502", x"500",
        x"4fe", x"4fc", x"4fa", x"4f8", x"4f6", x"4f4", x"4f2", x"4f0",
        x"4ee", x"4ec", x"4ea", x"4e8", x"4e6", x"4e4", x"4e2", x"4e0",
        x"4de", x"4dc", x"4da", x"4d8", x"4d6", x"4d4", x"4d2", x"4d0",
        x"4ce", x"4cc", x"4ca", x"4c8", x"4c6", x"4c4", x"4c2", x"4c0",
        x"4be", x"4bc", x"4ba", x"4b8", x"4b6", x"4b4", x"4b2", x"4b0",
        x"4ae", x"4ac", x"4aa", x"4a8", x"4a6", x"4a4", x"4a2", x"4a0",
        x"49e", x"49c", x"49a", x"498", x"496", x"494", x"492", x"490",
        x"48e", x"48c", x"48a", x"488", x"486", x"484", x"482", x"480",
        x"47e", x"47c", x"47a", x"478", x"476", x"474", x"472", x"470",
        x"46e", x"46c", x"46a", x"468", x"466", x"464", x"462", x"460",
        x"45e", x"45c", x"45a", x"458", x"456", x"454", x"452", x"450",
        x"44e", x"44c", x"44a", x"448", x"446", x"444", x"442", x"440",
        x"43e", x"43c", x"43a", x"438", x"436", x"434", x"432", x"430",
        x"42e", x"42c", x"42a", x"428", x"426", x"424", x"422", x"420",
        x"41e", x"41c", x"41a", x"418", x"416", x"414", x"412", x"410",
        x"40e", x"40c", x"40a", x"408", x"406", x"404", x"402", x"400",
        x"3fe", x"3fc", x"3fa", x"3f8", x"3f6", x"3f4", x"3f2", x"3f0",
        x"3ee", x"3ec", x"3ea", x"3e8", x"3e6", x"3e4", x"3e2", x"3e0",
        x"3de", x"3dc", x"3da", x"3d8", x"3d6", x"3d4", x"3d2", x"3d0",
        x"3ce", x"3cc", x"3ca", x"3c8", x"3c6", x"3c4", x"3c2", x"3c0",
        x"3be", x"3bc", x"3ba", x"3b8", x"3b6", x"3b4", x"3b2", x"3b0",
        x"3ae", x"3ac", x"3aa", x"3a8", x"3a6", x"3a4", x"3a2", x"3a0",
        x"39e", x"39c", x"39a", x"398", x"396", x"394", x"392", x"390",
        x"38e", x"38c", x"38a", x"388", x"386", x"384", x"382", x"380",
        x"37e", x"37c", x"37a", x"378", x"376", x"374", x"372", x"370",
        x"36e", x"36c", x"36a", x"368", x"366", x"364", x"362", x"360",
        x"35e", x"35c", x"35a", x"358", x"356", x"354", x"352", x"350",
        x"34e", x"34c", x"34a", x"348", x"346", x"344", x"342", x"340",
        x"33e", x"33c", x"33a", x"338", x"336", x"334", x"332", x"330",
        x"32e", x"32c", x"32a", x"328", x"326", x"324", x"322", x"320",
        x"31e", x"31c", x"31a", x"318", x"316", x"314", x"312", x"310",
        x"30e", x"30c", x"30a", x"308", x"306", x"304", x"302", x"300",
        x"2fe", x"2fc", x"2fa", x"2f8", x"2f6", x"2f4", x"2f2", x"2f0",
        x"2ee", x"2ec", x"2ea", x"2e8", x"2e6", x"2e4", x"2e2", x"2e0",
        x"2de", x"2dc", x"2da", x"2d8", x"2d6", x"2d4", x"2d2", x"2d0",
        x"2ce", x"2cc", x"2ca", x"2c8", x"2c6", x"2c4", x"2c2", x"2c0",
        x"2be", x"2bc", x"2ba", x"2b8", x"2b6", x"2b4", x"2b2", x"2b0",
        x"2ae", x"2ac", x"2aa", x"2a8", x"2a6", x"2a4", x"2a2", x"2a0",
        x"29e", x"29c", x"29a", x"298", x"296", x"294", x"292", x"290",
        x"28e", x"28c", x"28a", x"288", x"286", x"284", x"282", x"280",
        x"27e", x"27c", x"27a", x"278", x"276", x"274", x"272", x"270",
        x"26e", x"26c", x"26a", x"268", x"266", x"264", x"262", x"260",
        x"25e", x"25c", x"25a", x"258", x"256", x"254", x"252", x"250",
        x"24e", x"24c", x"24a", x"248", x"246", x"244", x"242", x"240",
        x"23e", x"23c", x"23a", x"238", x"236", x"234", x"232", x"230",
        x"22e", x"22c", x"22a", x"228", x"226", x"224", x"222", x"220",
        x"21e", x"21c", x"21a", x"218", x"216", x"214", x"212", x"210",
        x"20e", x"20c", x"20a", x"208", x"206", x"204", x"202", x"200",
        x"1fe", x"1fc", x"1fa", x"1f8", x"1f6", x"1f4", x"1f2", x"1f0",
        x"1ee", x"1ec", x"1ea", x"1e8", x"1e6", x"1e4", x"1e2", x"1e0",
        x"1de", x"1dc", x"1da", x"1d8", x"1d6", x"1d4", x"1d2", x"1d0",
        x"1ce", x"1cc", x"1ca", x"1c8", x"1c6", x"1c4", x"1c2", x"1c0",
        x"1be", x"1bc", x"1ba", x"1b8", x"1b6", x"1b4", x"1b2", x"1b0",
        x"1ae", x"1ac", x"1aa", x"1a8", x"1a6", x"1a4", x"1a2", x"1a0",
        x"19e", x"19c", x"19a", x"198", x"196", x"194", x"192", x"190",
        x"18e", x"18c", x"18a", x"188", x"186", x"184", x"182", x"180",
        x"17e", x"17c", x"17a", x"178", x"176", x"174", x"172", x"170",
        x"16e", x"16c", x"16a", x"168", x"166", x"164", x"162", x"160",
        x"15e", x"15c", x"15a", x"158", x"156", x"154", x"152", x"150",
        x"14e", x"14c", x"14a", x"148", x"146", x"144", x"142", x"140",
        x"13e", x"13c", x"13a", x"138", x"136", x"134", x"132", x"130",
        x"12e", x"12c", x"12a", x"128", x"126", x"124", x"122", x"120",
        x"11e", x"11c", x"11a", x"118", x"116", x"114", x"112", x"110",
        x"10e", x"10c", x"10a", x"108", x"106", x"104", x"102", x"100",
        x"0fe", x"0fc", x"0fa", x"0f8", x"0f6", x"0f4", x"0f2", x"0f0",
        x"0ee", x"0ec", x"0ea", x"0e8", x"0e6", x"0e4", x"0e2", x"0e0",
        x"0de", x"0dc", x"0da", x"0d8", x"0d6", x"0d4", x"0d2", x"0d0",
        x"0ce", x"0cc", x"0ca", x"0c8", x"0c6", x"0c4", x"0c2", x"0c0",
        x"0be", x"0bc", x"0ba", x"0b8", x"0b6", x"0b4", x"0b2", x"0b0",
        x"0ae", x"0ac", x"0aa", x"0a8", x"0a6", x"0a4", x"0a2", x"0a0",
        x"09e", x"09c", x"09a", x"098", x"096", x"094", x"092", x"090",
        x"08e", x"08c", x"08a", x"088", x"086", x"084", x"082", x"080",
        x"07e", x"07c", x"07a", x"078", x"076", x"074", x"072", x"070",
        x"06e", x"06c", x"06a", x"068", x"066", x"064", x"062", x"060",
        x"05e", x"05c", x"05a", x"058", x"056", x"054", x"052", x"050",
        x"04e", x"04c", x"04a", x"048", x"046", x"044", x"042", x"040",
        x"03e", x"03c", x"03a", x"038", x"036", x"034", x"032", x"030",
        x"02e", x"02c", x"02a", x"028", x"026", x"024", x"022", x"020",
        x"01e", x"01c", x"01a", x"018", x"016", x"014", x"012", x"010",
        x"00e", x"00c", x"00a", x"008", x"006", x"004", x"002", x"000"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr, clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp, en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
