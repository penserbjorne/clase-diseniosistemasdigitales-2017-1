library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom_triangulo is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(10 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom_triangulo;

architecture arch of rom_triangulo is
    type memoria_rom is array (0 to 2047) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"004", x"008", x"00c", x"010", x"014", x"018", x"01c", x"020",
        x"024", x"028", x"02c", x"030", x"034", x"038", x"03c", x"040",
        x"044", x"048", x"04c", x"050", x"054", x"058", x"05c", x"060",
        x"064", x"068", x"06c", x"070", x"074", x"078", x"07c", x"080",
        x"084", x"088", x"08c", x"090", x"094", x"098", x"09c", x"0a0",
        x"0a4", x"0a8", x"0ac", x"0b0", x"0b4", x"0b8", x"0bc", x"0c0",
        x"0c4", x"0c8", x"0cc", x"0d0", x"0d4", x"0d8", x"0dc", x"0e0",
        x"0e4", x"0e8", x"0ec", x"0f0", x"0f4", x"0f8", x"0fc", x"100",
        x"104", x"108", x"10c", x"110", x"114", x"118", x"11c", x"120",
        x"124", x"128", x"12c", x"130", x"134", x"138", x"13c", x"140",
        x"144", x"148", x"14c", x"150", x"154", x"158", x"15c", x"160",
        x"164", x"168", x"16c", x"170", x"174", x"178", x"17c", x"180",
        x"184", x"188", x"18c", x"190", x"194", x"198", x"19c", x"1a0",
        x"1a4", x"1a8", x"1ac", x"1b0", x"1b4", x"1b8", x"1bc", x"1c0",
        x"1c4", x"1c8", x"1cc", x"1d0", x"1d4", x"1d8", x"1dc", x"1e0",
        x"1e4", x"1e8", x"1ec", x"1f0", x"1f4", x"1f8", x"1fc", x"200",
        x"204", x"208", x"20c", x"210", x"214", x"218", x"21c", x"220",
        x"224", x"228", x"22c", x"230", x"234", x"238", x"23c", x"240",
        x"244", x"248", x"24c", x"250", x"254", x"258", x"25c", x"260",
        x"264", x"268", x"26c", x"270", x"274", x"278", x"27c", x"280",
        x"284", x"288", x"28c", x"290", x"294", x"298", x"29c", x"2a0",
        x"2a4", x"2a8", x"2ac", x"2b0", x"2b4", x"2b8", x"2bc", x"2c0",
        x"2c4", x"2c8", x"2cc", x"2d0", x"2d4", x"2d8", x"2dc", x"2e0",
        x"2e4", x"2e8", x"2ec", x"2f0", x"2f4", x"2f8", x"2fc", x"300",
        x"304", x"308", x"30c", x"310", x"314", x"318", x"31c", x"320",
        x"324", x"328", x"32c", x"330", x"334", x"338", x"33c", x"340",
        x"344", x"348", x"34c", x"350", x"354", x"358", x"35c", x"360",
        x"364", x"368", x"36c", x"370", x"374", x"378", x"37c", x"380",
        x"384", x"388", x"38c", x"390", x"394", x"398", x"39c", x"3a0",
        x"3a4", x"3a8", x"3ac", x"3b0", x"3b4", x"3b8", x"3bc", x"3c0",
        x"3c4", x"3c8", x"3cc", x"3d0", x"3d4", x"3d8", x"3dc", x"3e0",
        x"3e4", x"3e8", x"3ec", x"3f0", x"3f4", x"3f8", x"3fc", x"400",
        x"404", x"408", x"40c", x"410", x"414", x"418", x"41c", x"420",
        x"424", x"428", x"42c", x"430", x"434", x"438", x"43c", x"440",
        x"444", x"448", x"44c", x"450", x"454", x"458", x"45c", x"460",
        x"464", x"468", x"46c", x"470", x"474", x"478", x"47c", x"480",
        x"484", x"488", x"48c", x"490", x"494", x"498", x"49c", x"4a0",
        x"4a4", x"4a8", x"4ac", x"4b0", x"4b4", x"4b8", x"4bc", x"4c0",
        x"4c4", x"4c8", x"4cc", x"4d0", x"4d4", x"4d8", x"4dc", x"4e0",
        x"4e4", x"4e8", x"4ec", x"4f0", x"4f4", x"4f8", x"4fc", x"500",
        x"504", x"508", x"50c", x"510", x"514", x"518", x"51c", x"520",
        x"524", x"528", x"52c", x"530", x"534", x"538", x"53c", x"540",
        x"544", x"548", x"54c", x"550", x"554", x"558", x"55c", x"560",
        x"564", x"568", x"56c", x"570", x"574", x"578", x"57c", x"580",
        x"584", x"588", x"58c", x"590", x"594", x"598", x"59c", x"5a0",
        x"5a4", x"5a8", x"5ac", x"5b0", x"5b4", x"5b8", x"5bc", x"5c0",
        x"5c4", x"5c8", x"5cc", x"5d0", x"5d4", x"5d8", x"5dc", x"5e0",
        x"5e4", x"5e8", x"5ec", x"5f0", x"5f4", x"5f8", x"5fc", x"600",
        x"604", x"608", x"60c", x"610", x"614", x"618", x"61c", x"620",
        x"624", x"628", x"62c", x"630", x"634", x"638", x"63c", x"640",
        x"644", x"648", x"64c", x"650", x"654", x"658", x"65c", x"660",
        x"664", x"668", x"66c", x"670", x"674", x"678", x"67c", x"680",
        x"684", x"688", x"68c", x"690", x"694", x"698", x"69c", x"6a0",
        x"6a4", x"6a8", x"6ac", x"6b0", x"6b4", x"6b8", x"6bc", x"6c0",
        x"6c4", x"6c8", x"6cc", x"6d0", x"6d4", x"6d8", x"6dc", x"6e0",
        x"6e4", x"6e8", x"6ec", x"6f0", x"6f4", x"6f8", x"6fc", x"700",
        x"704", x"708", x"70c", x"710", x"714", x"718", x"71c", x"720",
        x"724", x"728", x"72c", x"730", x"734", x"738", x"73c", x"740",
        x"744", x"748", x"74c", x"750", x"754", x"758", x"75c", x"760",
        x"764", x"768", x"76c", x"770", x"774", x"778", x"77c", x"780",
        x"784", x"788", x"78c", x"790", x"794", x"798", x"79c", x"7a0",
        x"7a4", x"7a8", x"7ac", x"7b0", x"7b4", x"7b8", x"7bc", x"7c0",
        x"7c4", x"7c8", x"7cc", x"7d0", x"7d4", x"7d8", x"7dc", x"7e0",
        x"7e4", x"7e8", x"7ec", x"7f0", x"7f4", x"7f8", x"7fc", x"801",
        x"805", x"809", x"80d", x"811", x"815", x"819", x"81d", x"821",
        x"825", x"829", x"82d", x"831", x"835", x"839", x"83d", x"841",
        x"845", x"849", x"84d", x"851", x"855", x"859", x"85d", x"861",
        x"865", x"869", x"86d", x"871", x"875", x"879", x"87d", x"881",
        x"885", x"889", x"88d", x"891", x"895", x"899", x"89d", x"8a1",
        x"8a5", x"8a9", x"8ad", x"8b1", x"8b5", x"8b9", x"8bd", x"8c1",
        x"8c5", x"8c9", x"8cd", x"8d1", x"8d5", x"8d9", x"8dd", x"8e1",
        x"8e5", x"8e9", x"8ed", x"8f1", x"8f5", x"8f9", x"8fd", x"901",
        x"905", x"909", x"90d", x"911", x"915", x"919", x"91d", x"921",
        x"925", x"929", x"92d", x"931", x"935", x"939", x"93d", x"941",
        x"945", x"949", x"94d", x"951", x"955", x"959", x"95d", x"961",
        x"965", x"969", x"96d", x"971", x"975", x"979", x"97d", x"981",
        x"985", x"989", x"98d", x"991", x"995", x"999", x"99d", x"9a1",
        x"9a5", x"9a9", x"9ad", x"9b1", x"9b5", x"9b9", x"9bd", x"9c1",
        x"9c5", x"9c9", x"9cd", x"9d1", x"9d5", x"9d9", x"9dd", x"9e1",
        x"9e5", x"9e9", x"9ed", x"9f1", x"9f5", x"9f9", x"9fd", x"a01",
        x"a05", x"a09", x"a0d", x"a11", x"a15", x"a19", x"a1d", x"a21",
        x"a25", x"a29", x"a2d", x"a31", x"a35", x"a39", x"a3d", x"a41",
        x"a45", x"a49", x"a4d", x"a51", x"a55", x"a59", x"a5d", x"a61",
        x"a65", x"a69", x"a6d", x"a71", x"a75", x"a79", x"a7d", x"a81",
        x"a85", x"a89", x"a8d", x"a91", x"a95", x"a99", x"a9d", x"aa1",
        x"aa5", x"aa9", x"aad", x"ab1", x"ab5", x"ab9", x"abd", x"ac1",
        x"ac5", x"ac9", x"acd", x"ad1", x"ad5", x"ad9", x"add", x"ae1",
        x"ae5", x"ae9", x"aed", x"af1", x"af5", x"af9", x"afd", x"b01",
        x"b05", x"b09", x"b0d", x"b11", x"b15", x"b19", x"b1d", x"b21",
        x"b25", x"b29", x"b2d", x"b31", x"b35", x"b39", x"b3d", x"b41",
        x"b45", x"b49", x"b4d", x"b51", x"b55", x"b59", x"b5d", x"b61",
        x"b65", x"b69", x"b6d", x"b71", x"b75", x"b79", x"b7d", x"b81",
        x"b85", x"b89", x"b8d", x"b91", x"b95", x"b99", x"b9d", x"ba1",
        x"ba5", x"ba9", x"bad", x"bb1", x"bb5", x"bb9", x"bbd", x"bc1",
        x"bc5", x"bc9", x"bcd", x"bd1", x"bd5", x"bd9", x"bdd", x"be1",
        x"be5", x"be9", x"bed", x"bf1", x"bf5", x"bf9", x"bfd", x"c01",
        x"c05", x"c09", x"c0d", x"c11", x"c15", x"c19", x"c1d", x"c21",
        x"c25", x"c29", x"c2d", x"c31", x"c35", x"c39", x"c3d", x"c41",
        x"c45", x"c49", x"c4d", x"c51", x"c55", x"c59", x"c5d", x"c61",
        x"c65", x"c69", x"c6d", x"c71", x"c75", x"c79", x"c7d", x"c81",
        x"c85", x"c89", x"c8d", x"c91", x"c95", x"c99", x"c9d", x"ca1",
        x"ca5", x"ca9", x"cad", x"cb1", x"cb5", x"cb9", x"cbd", x"cc1",
        x"cc5", x"cc9", x"ccd", x"cd1", x"cd5", x"cd9", x"cdd", x"ce1",
        x"ce5", x"ce9", x"ced", x"cf1", x"cf5", x"cf9", x"cfd", x"d01",
        x"d05", x"d09", x"d0d", x"d11", x"d15", x"d19", x"d1d", x"d21",
        x"d25", x"d29", x"d2d", x"d31", x"d35", x"d39", x"d3d", x"d41",
        x"d45", x"d49", x"d4d", x"d51", x"d55", x"d59", x"d5d", x"d61",
        x"d65", x"d69", x"d6d", x"d71", x"d75", x"d79", x"d7d", x"d81",
        x"d85", x"d89", x"d8d", x"d91", x"d95", x"d99", x"d9d", x"da1",
        x"da5", x"da9", x"dad", x"db1", x"db5", x"db9", x"dbd", x"dc1",
        x"dc5", x"dc9", x"dcd", x"dd1", x"dd5", x"dd9", x"ddd", x"de1",
        x"de5", x"de9", x"ded", x"df1", x"df5", x"df9", x"dfd", x"e01",
        x"e05", x"e09", x"e0d", x"e11", x"e15", x"e19", x"e1d", x"e21",
        x"e25", x"e29", x"e2d", x"e31", x"e35", x"e39", x"e3d", x"e41",
        x"e45", x"e49", x"e4d", x"e51", x"e55", x"e59", x"e5d", x"e61",
        x"e65", x"e69", x"e6d", x"e71", x"e75", x"e79", x"e7d", x"e81",
        x"e85", x"e89", x"e8d", x"e91", x"e95", x"e99", x"e9d", x"ea1",
        x"ea5", x"ea9", x"ead", x"eb1", x"eb5", x"eb9", x"ebd", x"ec1",
        x"ec5", x"ec9", x"ecd", x"ed1", x"ed5", x"ed9", x"edd", x"ee1",
        x"ee5", x"ee9", x"eed", x"ef1", x"ef5", x"ef9", x"efd", x"f01",
        x"f05", x"f09", x"f0d", x"f11", x"f15", x"f19", x"f1d", x"f21",
        x"f25", x"f29", x"f2d", x"f31", x"f35", x"f39", x"f3d", x"f41",
        x"f45", x"f49", x"f4d", x"f51", x"f55", x"f59", x"f5d", x"f61",
        x"f65", x"f69", x"f6d", x"f71", x"f75", x"f79", x"f7d", x"f81",
        x"f85", x"f89", x"f8d", x"f91", x"f95", x"f99", x"f9d", x"fa1",
        x"fa5", x"fa9", x"fad", x"fb1", x"fb5", x"fb9", x"fbd", x"fc1",
        x"fc5", x"fc9", x"fcd", x"fd1", x"fd5", x"fd9", x"fdd", x"fe1",
        x"fe5", x"fe9", x"fed", x"ff1", x"ff5", x"ff9", x"ffd", x"fff",
        x"ffd", x"ff9", x"ff5", x"ff1", x"fed", x"fe9", x"fe5", x"fe1",
        x"fdd", x"fd9", x"fd5", x"fd1", x"fcd", x"fc9", x"fc5", x"fc1",
        x"fbd", x"fb9", x"fb5", x"fb1", x"fad", x"fa9", x"fa5", x"fa1",
        x"f9d", x"f99", x"f95", x"f91", x"f8d", x"f89", x"f85", x"f81",
        x"f7d", x"f79", x"f75", x"f71", x"f6d", x"f69", x"f65", x"f61",
        x"f5d", x"f59", x"f55", x"f51", x"f4d", x"f49", x"f45", x"f41",
        x"f3d", x"f39", x"f35", x"f31", x"f2d", x"f29", x"f25", x"f21",
        x"f1d", x"f19", x"f15", x"f11", x"f0d", x"f09", x"f05", x"f01",
        x"efd", x"ef9", x"ef5", x"ef1", x"eed", x"ee9", x"ee5", x"ee1",
        x"edd", x"ed9", x"ed5", x"ed1", x"ecd", x"ec9", x"ec5", x"ec1",
        x"ebd", x"eb9", x"eb5", x"eb1", x"ead", x"ea9", x"ea5", x"ea1",
        x"e9d", x"e99", x"e95", x"e91", x"e8d", x"e89", x"e85", x"e81",
        x"e7d", x"e79", x"e75", x"e71", x"e6d", x"e69", x"e65", x"e61",
        x"e5d", x"e59", x"e55", x"e51", x"e4d", x"e49", x"e45", x"e41",
        x"e3d", x"e39", x"e35", x"e31", x"e2d", x"e29", x"e25", x"e21",
        x"e1d", x"e19", x"e15", x"e11", x"e0d", x"e09", x"e05", x"e01",
        x"dfd", x"df9", x"df5", x"df1", x"ded", x"de9", x"de5", x"de1",
        x"ddd", x"dd9", x"dd5", x"dd1", x"dcd", x"dc9", x"dc5", x"dc1",
        x"dbd", x"db9", x"db5", x"db1", x"dad", x"da9", x"da5", x"da1",
        x"d9d", x"d99", x"d95", x"d91", x"d8d", x"d89", x"d85", x"d81",
        x"d7d", x"d79", x"d75", x"d71", x"d6d", x"d69", x"d65", x"d61",
        x"d5d", x"d59", x"d55", x"d51", x"d4d", x"d49", x"d45", x"d41",
        x"d3d", x"d39", x"d35", x"d31", x"d2d", x"d29", x"d25", x"d21",
        x"d1d", x"d19", x"d15", x"d11", x"d0d", x"d09", x"d05", x"d01",
        x"cfd", x"cf9", x"cf5", x"cf1", x"ced", x"ce9", x"ce5", x"ce1",
        x"cdd", x"cd9", x"cd5", x"cd1", x"ccd", x"cc9", x"cc5", x"cc1",
        x"cbd", x"cb9", x"cb5", x"cb1", x"cad", x"ca9", x"ca5", x"ca1",
        x"c9d", x"c99", x"c95", x"c91", x"c8d", x"c89", x"c85", x"c81",
        x"c7d", x"c79", x"c75", x"c71", x"c6d", x"c69", x"c65", x"c61",
        x"c5d", x"c59", x"c55", x"c51", x"c4d", x"c49", x"c45", x"c41",
        x"c3d", x"c39", x"c35", x"c31", x"c2d", x"c29", x"c25", x"c21",
        x"c1d", x"c19", x"c15", x"c11", x"c0d", x"c09", x"c05", x"c01",
        x"bfd", x"bf9", x"bf5", x"bf1", x"bed", x"be9", x"be5", x"be1",
        x"bdd", x"bd9", x"bd5", x"bd1", x"bcd", x"bc9", x"bc5", x"bc1",
        x"bbd", x"bb9", x"bb5", x"bb1", x"bad", x"ba9", x"ba5", x"ba1",
        x"b9d", x"b99", x"b95", x"b91", x"b8d", x"b89", x"b85", x"b81",
        x"b7d", x"b79", x"b75", x"b71", x"b6d", x"b69", x"b65", x"b61",
        x"b5d", x"b59", x"b55", x"b51", x"b4d", x"b49", x"b45", x"b41",
        x"b3d", x"b39", x"b35", x"b31", x"b2d", x"b29", x"b25", x"b21",
        x"b1d", x"b19", x"b15", x"b11", x"b0d", x"b09", x"b05", x"b01",
        x"afd", x"af9", x"af5", x"af1", x"aed", x"ae9", x"ae5", x"ae1",
        x"add", x"ad9", x"ad5", x"ad1", x"acd", x"ac9", x"ac5", x"ac1",
        x"abd", x"ab9", x"ab5", x"ab1", x"aad", x"aa9", x"aa5", x"aa1",
        x"a9d", x"a99", x"a95", x"a91", x"a8d", x"a89", x"a85", x"a81",
        x"a7d", x"a79", x"a75", x"a71", x"a6d", x"a69", x"a65", x"a61",
        x"a5d", x"a59", x"a55", x"a51", x"a4d", x"a49", x"a45", x"a41",
        x"a3d", x"a39", x"a35", x"a31", x"a2d", x"a29", x"a25", x"a21",
        x"a1d", x"a19", x"a15", x"a11", x"a0d", x"a09", x"a05", x"a01",
        x"9fd", x"9f9", x"9f5", x"9f1", x"9ed", x"9e9", x"9e5", x"9e1",
        x"9dd", x"9d9", x"9d5", x"9d1", x"9cd", x"9c9", x"9c5", x"9c1",
        x"9bd", x"9b9", x"9b5", x"9b1", x"9ad", x"9a9", x"9a5", x"9a1",
        x"99d", x"999", x"995", x"991", x"98d", x"989", x"985", x"981",
        x"97d", x"979", x"975", x"971", x"96d", x"969", x"965", x"961",
        x"95d", x"959", x"955", x"951", x"94d", x"949", x"945", x"941",
        x"93d", x"939", x"935", x"931", x"92d", x"929", x"925", x"921",
        x"91d", x"919", x"915", x"911", x"90d", x"909", x"905", x"901",
        x"8fd", x"8f9", x"8f5", x"8f1", x"8ed", x"8e9", x"8e5", x"8e1",
        x"8dd", x"8d9", x"8d5", x"8d1", x"8cd", x"8c9", x"8c5", x"8c1",
        x"8bd", x"8b9", x"8b5", x"8b1", x"8ad", x"8a9", x"8a5", x"8a1",
        x"89d", x"899", x"895", x"891", x"88d", x"889", x"885", x"881",
        x"87d", x"879", x"875", x"871", x"86d", x"869", x"865", x"861",
        x"85d", x"859", x"855", x"851", x"84d", x"849", x"845", x"841",
        x"83d", x"839", x"835", x"831", x"82d", x"829", x"825", x"821",
        x"81d", x"819", x"815", x"811", x"80d", x"809", x"805", x"801",
        x"7fc", x"7f8", x"7f4", x"7f0", x"7ec", x"7e8", x"7e4", x"7e0",
        x"7dc", x"7d8", x"7d4", x"7d0", x"7cc", x"7c8", x"7c4", x"7c0",
        x"7bc", x"7b8", x"7b4", x"7b0", x"7ac", x"7a8", x"7a4", x"7a0",
        x"79c", x"798", x"794", x"790", x"78c", x"788", x"784", x"780",
        x"77c", x"778", x"774", x"770", x"76c", x"768", x"764", x"760",
        x"75c", x"758", x"754", x"750", x"74c", x"748", x"744", x"740",
        x"73c", x"738", x"734", x"730", x"72c", x"728", x"724", x"720",
        x"71c", x"718", x"714", x"710", x"70c", x"708", x"704", x"700",
        x"6fc", x"6f8", x"6f4", x"6f0", x"6ec", x"6e8", x"6e4", x"6e0",
        x"6dc", x"6d8", x"6d4", x"6d0", x"6cc", x"6c8", x"6c4", x"6c0",
        x"6bc", x"6b8", x"6b4", x"6b0", x"6ac", x"6a8", x"6a4", x"6a0",
        x"69c", x"698", x"694", x"690", x"68c", x"688", x"684", x"680",
        x"67c", x"678", x"674", x"670", x"66c", x"668", x"664", x"660",
        x"65c", x"658", x"654", x"650", x"64c", x"648", x"644", x"640",
        x"63c", x"638", x"634", x"630", x"62c", x"628", x"624", x"620",
        x"61c", x"618", x"614", x"610", x"60c", x"608", x"604", x"600",
        x"5fc", x"5f8", x"5f4", x"5f0", x"5ec", x"5e8", x"5e4", x"5e0",
        x"5dc", x"5d8", x"5d4", x"5d0", x"5cc", x"5c8", x"5c4", x"5c0",
        x"5bc", x"5b8", x"5b4", x"5b0", x"5ac", x"5a8", x"5a4", x"5a0",
        x"59c", x"598", x"594", x"590", x"58c", x"588", x"584", x"580",
        x"57c", x"578", x"574", x"570", x"56c", x"568", x"564", x"560",
        x"55c", x"558", x"554", x"550", x"54c", x"548", x"544", x"540",
        x"53c", x"538", x"534", x"530", x"52c", x"528", x"524", x"520",
        x"51c", x"518", x"514", x"510", x"50c", x"508", x"504", x"500",
        x"4fc", x"4f8", x"4f4", x"4f0", x"4ec", x"4e8", x"4e4", x"4e0",
        x"4dc", x"4d8", x"4d4", x"4d0", x"4cc", x"4c8", x"4c4", x"4c0",
        x"4bc", x"4b8", x"4b4", x"4b0", x"4ac", x"4a8", x"4a4", x"4a0",
        x"49c", x"498", x"494", x"490", x"48c", x"488", x"484", x"480",
        x"47c", x"478", x"474", x"470", x"46c", x"468", x"464", x"460",
        x"45c", x"458", x"454", x"450", x"44c", x"448", x"444", x"440",
        x"43c", x"438", x"434", x"430", x"42c", x"428", x"424", x"420",
        x"41c", x"418", x"414", x"410", x"40c", x"408", x"404", x"400",
        x"3fc", x"3f8", x"3f4", x"3f0", x"3ec", x"3e8", x"3e4", x"3e0",
        x"3dc", x"3d8", x"3d4", x"3d0", x"3cc", x"3c8", x"3c4", x"3c0",
        x"3bc", x"3b8", x"3b4", x"3b0", x"3ac", x"3a8", x"3a4", x"3a0",
        x"39c", x"398", x"394", x"390", x"38c", x"388", x"384", x"380",
        x"37c", x"378", x"374", x"370", x"36c", x"368", x"364", x"360",
        x"35c", x"358", x"354", x"350", x"34c", x"348", x"344", x"340",
        x"33c", x"338", x"334", x"330", x"32c", x"328", x"324", x"320",
        x"31c", x"318", x"314", x"310", x"30c", x"308", x"304", x"300",
        x"2fc", x"2f8", x"2f4", x"2f0", x"2ec", x"2e8", x"2e4", x"2e0",
        x"2dc", x"2d8", x"2d4", x"2d0", x"2cc", x"2c8", x"2c4", x"2c0",
        x"2bc", x"2b8", x"2b4", x"2b0", x"2ac", x"2a8", x"2a4", x"2a0",
        x"29c", x"298", x"294", x"290", x"28c", x"288", x"284", x"280",
        x"27c", x"278", x"274", x"270", x"26c", x"268", x"264", x"260",
        x"25c", x"258", x"254", x"250", x"24c", x"248", x"244", x"240",
        x"23c", x"238", x"234", x"230", x"22c", x"228", x"224", x"220",
        x"21c", x"218", x"214", x"210", x"20c", x"208", x"204", x"200",
        x"1fc", x"1f8", x"1f4", x"1f0", x"1ec", x"1e8", x"1e4", x"1e0",
        x"1dc", x"1d8", x"1d4", x"1d0", x"1cc", x"1c8", x"1c4", x"1c0",
        x"1bc", x"1b8", x"1b4", x"1b0", x"1ac", x"1a8", x"1a4", x"1a0",
        x"19c", x"198", x"194", x"190", x"18c", x"188", x"184", x"180",
        x"17c", x"178", x"174", x"170", x"16c", x"168", x"164", x"160",
        x"15c", x"158", x"154", x"150", x"14c", x"148", x"144", x"140",
        x"13c", x"138", x"134", x"130", x"12c", x"128", x"124", x"120",
        x"11c", x"118", x"114", x"110", x"10c", x"108", x"104", x"100",
        x"0fc", x"0f8", x"0f4", x"0f0", x"0ec", x"0e8", x"0e4", x"0e0",
        x"0dc", x"0d8", x"0d4", x"0d0", x"0cc", x"0c8", x"0c4", x"0c0",
        x"0bc", x"0b8", x"0b4", x"0b0", x"0ac", x"0a8", x"0a4", x"0a0",
        x"09c", x"098", x"094", x"090", x"08c", x"088", x"084", x"080",
        x"07c", x"078", x"074", x"070", x"06c", x"068", x"064", x"060",
        x"05c", x"058", x"054", x"050", x"04c", x"048", x"044", x"040",
        x"03c", x"038", x"034", x"030", x"02c", x"028", x"024", x"020",
        x"01c", x"018", x"014", x"010", x"00c", x"008", x"004", x"000"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr, clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp, en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
