library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(10 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom;

architecture arch of rom is
    type memoria_rom is array (0 to 2047) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"001", x"002", x"003", x"004", x"005", x"006", x"007", x"008",
        x"009", x"00a", x"00b", x"00c", x"00d", x"00e", x"00f", x"010",
        x"011", x"012", x"013", x"014", x"015", x"016", x"017", x"018",
        x"019", x"01a", x"01b", x"01c", x"01d", x"01e", x"01f", x"020",
        x"021", x"022", x"023", x"024", x"025", x"026", x"027", x"028",
        x"029", x"02a", x"02b", x"02c", x"02d", x"02e", x"02f", x"030",
        x"031", x"032", x"033", x"034", x"035", x"036", x"037", x"038",
        x"039", x"03a", x"03b", x"03c", x"03d", x"03e", x"03f", x"040",
        x"041", x"042", x"043", x"044", x"045", x"046", x"047", x"048",
        x"049", x"04a", x"04b", x"04c", x"04d", x"04e", x"04f", x"050",
        x"051", x"052", x"053", x"054", x"055", x"056", x"057", x"058",
        x"059", x"05a", x"05b", x"05c", x"05d", x"05e", x"05f", x"060",
        x"061", x"062", x"063", x"064", x"065", x"066", x"067", x"068",
        x"069", x"06a", x"06b", x"06c", x"06d", x"06e", x"06f", x"070",
        x"071", x"072", x"073", x"074", x"075", x"076", x"077", x"078",
        x"079", x"07a", x"07b", x"07c", x"07d", x"07e", x"07f", x"080",
        x"081", x"082", x"083", x"084", x"085", x"086", x"087", x"088",
        x"089", x"08a", x"08b", x"08c", x"08d", x"08e", x"08f", x"090",
        x"091", x"092", x"093", x"094", x"095", x"096", x"097", x"098",
        x"099", x"09a", x"09b", x"09c", x"09d", x"09e", x"09f", x"0a0",
        x"0a1", x"0a2", x"0a3", x"0a4", x"0a5", x"0a6", x"0a7", x"0a8",
        x"0a9", x"0aa", x"0ab", x"0ac", x"0ad", x"0ae", x"0af", x"0b0",
        x"0b1", x"0b2", x"0b3", x"0b4", x"0b5", x"0b6", x"0b7", x"0b8",
        x"0b9", x"0ba", x"0bb", x"0bc", x"0bd", x"0be", x"0bf", x"0c0",
        x"0c1", x"0c2", x"0c3", x"0c4", x"0c5", x"0c6", x"0c7", x"0c8",
        x"0c9", x"0ca", x"0cb", x"0cc", x"0cd", x"0ce", x"0cf", x"0d0",
        x"0d1", x"0d2", x"0d3", x"0d4", x"0d5", x"0d6", x"0d7", x"0d8",
        x"0d9", x"0da", x"0db", x"0dc", x"0dd", x"0de", x"0df", x"0e0",
        x"0e1", x"0e2", x"0e3", x"0e4", x"0e5", x"0e6", x"0e7", x"0e8",
        x"0e9", x"0ea", x"0eb", x"0ec", x"0ed", x"0ee", x"0ef", x"0f0",
        x"0f1", x"0f2", x"0f3", x"0f4", x"0f5", x"0f6", x"0f7", x"0f8",
        x"0f9", x"0fa", x"0fb", x"0fc", x"0fd", x"0fe", x"0ff", x"100",
        x"101", x"102", x"103", x"104", x"105", x"106", x"107", x"108",
        x"109", x"10a", x"10b", x"10c", x"10d", x"10e", x"10f", x"110",
        x"111", x"112", x"113", x"114", x"115", x"116", x"117", x"118",
        x"119", x"11a", x"11b", x"11c", x"11d", x"11e", x"11f", x"120",
        x"121", x"122", x"123", x"124", x"125", x"126", x"127", x"128",
        x"129", x"12a", x"12b", x"12c", x"12d", x"12e", x"12f", x"130",
        x"131", x"132", x"133", x"134", x"135", x"136", x"137", x"138",
        x"139", x"13a", x"13b", x"13c", x"13d", x"13e", x"13f", x"140",
        x"141", x"142", x"143", x"144", x"145", x"146", x"147", x"148",
        x"149", x"14a", x"14b", x"14c", x"14d", x"14e", x"14f", x"150",
        x"151", x"152", x"153", x"154", x"155", x"156", x"157", x"158",
        x"159", x"15a", x"15b", x"15c", x"15d", x"15e", x"15f", x"160",
        x"161", x"162", x"163", x"164", x"165", x"166", x"167", x"168",
        x"169", x"16a", x"16b", x"16c", x"16d", x"16e", x"16f", x"170",
        x"171", x"172", x"173", x"174", x"175", x"176", x"177", x"178",
        x"179", x"17a", x"17b", x"17c", x"17d", x"17e", x"17f", x"180",
        x"181", x"182", x"183", x"184", x"185", x"186", x"187", x"188",
        x"189", x"18a", x"18b", x"18c", x"18d", x"18e", x"18f", x"190",
        x"191", x"192", x"193", x"194", x"195", x"196", x"197", x"198",
        x"199", x"19a", x"19b", x"19c", x"19d", x"19e", x"19f", x"1a0",
        x"1a1", x"1a2", x"1a3", x"1a4", x"1a5", x"1a6", x"1a7", x"1a8",
        x"1a9", x"1aa", x"1ab", x"1ac", x"1ad", x"1ae", x"1af", x"1b0",
        x"1b1", x"1b2", x"1b3", x"1b4", x"1b5", x"1b6", x"1b7", x"1b8",
        x"1b9", x"1ba", x"1bb", x"1bc", x"1bd", x"1be", x"1bf", x"1c0",
        x"1c1", x"1c2", x"1c3", x"1c4", x"1c5", x"1c6", x"1c7", x"1c8",
        x"1c9", x"1ca", x"1cb", x"1cc", x"1cd", x"1ce", x"1cf", x"1d0",
        x"1d1", x"1d2", x"1d3", x"1d4", x"1d5", x"1d6", x"1d7", x"1d8",
        x"1d9", x"1da", x"1db", x"1dc", x"1dd", x"1de", x"1df", x"1e0",
        x"1e1", x"1e2", x"1e3", x"1e4", x"1e5", x"1e6", x"1e7", x"1e8",
        x"1e9", x"1ea", x"1eb", x"1ec", x"1ed", x"1ee", x"1ef", x"1f0",
        x"1f1", x"1f2", x"1f3", x"1f4", x"1f5", x"1f6", x"1f7", x"1f8",
        x"1f9", x"1fa", x"1fb", x"1fc", x"1fd", x"1fe", x"1ff", x"200",
        x"201", x"202", x"203", x"204", x"205", x"206", x"207", x"208",
        x"209", x"20a", x"20b", x"20c", x"20d", x"20e", x"20f", x"210",
        x"211", x"212", x"213", x"214", x"215", x"216", x"217", x"218",
        x"219", x"21a", x"21b", x"21c", x"21d", x"21e", x"21f", x"220",
        x"221", x"222", x"223", x"224", x"225", x"226", x"227", x"228",
        x"229", x"22a", x"22b", x"22c", x"22d", x"22e", x"22f", x"230",
        x"231", x"232", x"233", x"234", x"235", x"236", x"237", x"238",
        x"239", x"23a", x"23b", x"23c", x"23d", x"23e", x"23f", x"240",
        x"241", x"242", x"243", x"244", x"245", x"246", x"247", x"248",
        x"249", x"24a", x"24b", x"24c", x"24d", x"24e", x"24f", x"250",
        x"251", x"252", x"253", x"254", x"255", x"256", x"257", x"258",
        x"259", x"25a", x"25b", x"25c", x"25d", x"25e", x"25f", x"260",
        x"261", x"262", x"263", x"264", x"265", x"266", x"267", x"268",
        x"269", x"26a", x"26b", x"26c", x"26d", x"26e", x"26f", x"270",
        x"271", x"272", x"273", x"274", x"275", x"276", x"277", x"278",
        x"279", x"27a", x"27b", x"27c", x"27d", x"27e", x"27f", x"280",
        x"281", x"282", x"283", x"284", x"285", x"286", x"287", x"288",
        x"289", x"28a", x"28b", x"28c", x"28d", x"28e", x"28f", x"290",
        x"291", x"292", x"293", x"294", x"295", x"296", x"297", x"298",
        x"299", x"29a", x"29b", x"29c", x"29d", x"29e", x"29f", x"2a0",
        x"2a1", x"2a2", x"2a3", x"2a4", x"2a5", x"2a6", x"2a7", x"2a8",
        x"2a9", x"2aa", x"2ab", x"2ac", x"2ad", x"2ae", x"2af", x"2b0",
        x"2b1", x"2b2", x"2b3", x"2b4", x"2b5", x"2b6", x"2b7", x"2b8",
        x"2b9", x"2ba", x"2bb", x"2bc", x"2bd", x"2be", x"2bf", x"2c0",
        x"2c1", x"2c2", x"2c3", x"2c4", x"2c5", x"2c6", x"2c7", x"2c8",
        x"2c9", x"2ca", x"2cb", x"2cc", x"2cd", x"2ce", x"2cf", x"2d0",
        x"2d1", x"2d2", x"2d3", x"2d4", x"2d5", x"2d6", x"2d7", x"2d8",
        x"2d9", x"2da", x"2db", x"2dc", x"2dd", x"2de", x"2df", x"2e0",
        x"2e1", x"2e2", x"2e3", x"2e4", x"2e5", x"2e6", x"2e7", x"2e8",
        x"2e9", x"2ea", x"2eb", x"2ec", x"2ed", x"2ee", x"2ef", x"2f0",
        x"2f1", x"2f2", x"2f3", x"2f4", x"2f5", x"2f6", x"2f7", x"2f8",
        x"2f9", x"2fa", x"2fb", x"2fc", x"2fd", x"2fe", x"2ff", x"300",
        x"301", x"302", x"303", x"304", x"305", x"306", x"307", x"308",
        x"309", x"30a", x"30b", x"30c", x"30d", x"30e", x"30f", x"310",
        x"311", x"312", x"313", x"314", x"315", x"316", x"317", x"318",
        x"319", x"31a", x"31b", x"31c", x"31d", x"31e", x"31f", x"320",
        x"321", x"322", x"323", x"324", x"325", x"326", x"327", x"328",
        x"329", x"32a", x"32b", x"32c", x"32d", x"32e", x"32f", x"330",
        x"331", x"332", x"333", x"334", x"335", x"336", x"337", x"338",
        x"339", x"33a", x"33b", x"33c", x"33d", x"33e", x"33f", x"340",
        x"341", x"342", x"343", x"344", x"345", x"346", x"347", x"348",
        x"349", x"34a", x"34b", x"34c", x"34d", x"34e", x"34f", x"350",
        x"351", x"352", x"353", x"354", x"355", x"356", x"357", x"358",
        x"359", x"35a", x"35b", x"35c", x"35d", x"35e", x"35f", x"360",
        x"361", x"362", x"363", x"364", x"365", x"366", x"367", x"368",
        x"369", x"36a", x"36b", x"36c", x"36d", x"36e", x"36f", x"370",
        x"371", x"372", x"373", x"374", x"375", x"376", x"377", x"378",
        x"379", x"37a", x"37b", x"37c", x"37d", x"37e", x"37f", x"380",
        x"381", x"382", x"383", x"384", x"385", x"386", x"387", x"388",
        x"389", x"38a", x"38b", x"38c", x"38d", x"38e", x"38f", x"390",
        x"391", x"392", x"393", x"394", x"395", x"396", x"397", x"398",
        x"399", x"39a", x"39b", x"39c", x"39d", x"39e", x"39f", x"3a0",
        x"3a1", x"3a2", x"3a3", x"3a4", x"3a5", x"3a6", x"3a7", x"3a8",
        x"3a9", x"3aa", x"3ab", x"3ac", x"3ad", x"3ae", x"3af", x"3b0",
        x"3b1", x"3b2", x"3b3", x"3b4", x"3b5", x"3b6", x"3b7", x"3b8",
        x"3b9", x"3ba", x"3bb", x"3bc", x"3bd", x"3be", x"3bf", x"3c0",
        x"3c1", x"3c2", x"3c3", x"3c4", x"3c5", x"3c6", x"3c7", x"3c8",
        x"3c9", x"3ca", x"3cb", x"3cc", x"3cd", x"3ce", x"3cf", x"3d0",
        x"3d1", x"3d2", x"3d3", x"3d4", x"3d5", x"3d6", x"3d7", x"3d8",
        x"3d9", x"3da", x"3db", x"3dc", x"3dd", x"3de", x"3df", x"3e0",
        x"3e1", x"3e2", x"3e3", x"3e4", x"3e5", x"3e6", x"3e7", x"3e8",
        x"3e9", x"3ea", x"3eb", x"3ec", x"3ed", x"3ee", x"3ef", x"3f0",
        x"3f1", x"3f2", x"3f3", x"3f4", x"3f5", x"3f6", x"3f7", x"3f8",
        x"3f9", x"3fa", x"3fb", x"3fc", x"3fd", x"3fe", x"3ff", x"400",
        x"401", x"402", x"403", x"404", x"405", x"406", x"407", x"408",
        x"409", x"40a", x"40b", x"40c", x"40d", x"40e", x"40f", x"410",
        x"411", x"412", x"413", x"414", x"415", x"416", x"417", x"418",
        x"419", x"41a", x"41b", x"41c", x"41d", x"41e", x"41f", x"420",
        x"421", x"422", x"423", x"424", x"425", x"426", x"427", x"428",
        x"429", x"42a", x"42b", x"42c", x"42d", x"42e", x"42f", x"430",
        x"431", x"432", x"433", x"434", x"435", x"436", x"437", x"438",
        x"439", x"43a", x"43b", x"43c", x"43d", x"43e", x"43f", x"440",
        x"441", x"442", x"443", x"444", x"445", x"446", x"447", x"448",
        x"449", x"44a", x"44b", x"44c", x"44d", x"44e", x"44f", x"450",
        x"451", x"452", x"453", x"454", x"455", x"456", x"457", x"458",
        x"459", x"45a", x"45b", x"45c", x"45d", x"45e", x"45f", x"460",
        x"461", x"462", x"463", x"464", x"465", x"466", x"467", x"468",
        x"469", x"46a", x"46b", x"46c", x"46d", x"46e", x"46f", x"470",
        x"471", x"472", x"473", x"474", x"475", x"476", x"477", x"478",
        x"479", x"47a", x"47b", x"47c", x"47d", x"47e", x"47f", x"480",
        x"481", x"482", x"483", x"484", x"485", x"486", x"487", x"488",
        x"489", x"48a", x"48b", x"48c", x"48d", x"48e", x"48f", x"490",
        x"491", x"492", x"493", x"494", x"495", x"496", x"497", x"498",
        x"499", x"49a", x"49b", x"49c", x"49d", x"49e", x"49f", x"4a0",
        x"4a1", x"4a2", x"4a3", x"4a4", x"4a5", x"4a6", x"4a7", x"4a8",
        x"4a9", x"4aa", x"4ab", x"4ac", x"4ad", x"4ae", x"4af", x"4b0",
        x"4b1", x"4b2", x"4b3", x"4b4", x"4b5", x"4b6", x"4b7", x"4b8",
        x"4b9", x"4ba", x"4bb", x"4bc", x"4bd", x"4be", x"4bf", x"4c0",
        x"4c1", x"4c2", x"4c3", x"4c4", x"4c5", x"4c6", x"4c7", x"4c8",
        x"4c9", x"4ca", x"4cb", x"4cc", x"4cd", x"4ce", x"4cf", x"4d0",
        x"4d1", x"4d2", x"4d3", x"4d4", x"4d5", x"4d6", x"4d7", x"4d8",
        x"4d9", x"4da", x"4db", x"4dc", x"4dd", x"4de", x"4df", x"4e0",
        x"4e1", x"4e2", x"4e3", x"4e4", x"4e5", x"4e6", x"4e7", x"4e8",
        x"4e9", x"4ea", x"4eb", x"4ec", x"4ed", x"4ee", x"4ef", x"4f0",
        x"4f1", x"4f2", x"4f3", x"4f4", x"4f5", x"4f6", x"4f7", x"4f8",
        x"4f9", x"4fa", x"4fb", x"4fc", x"4fd", x"4fe", x"4ff", x"500",
        x"501", x"502", x"503", x"504", x"505", x"506", x"507", x"508",
        x"509", x"50a", x"50b", x"50c", x"50d", x"50e", x"50f", x"510",
        x"511", x"512", x"513", x"514", x"515", x"516", x"517", x"518",
        x"519", x"51a", x"51b", x"51c", x"51d", x"51e", x"51f", x"520",
        x"521", x"522", x"523", x"524", x"525", x"526", x"527", x"528",
        x"529", x"52a", x"52b", x"52c", x"52d", x"52e", x"52f", x"530",
        x"531", x"532", x"533", x"534", x"535", x"536", x"537", x"538",
        x"539", x"53a", x"53b", x"53c", x"53d", x"53e", x"53f", x"540",
        x"541", x"542", x"543", x"544", x"545", x"546", x"547", x"548",
        x"549", x"54a", x"54b", x"54c", x"54d", x"54e", x"54f", x"550",
        x"551", x"552", x"553", x"554", x"555", x"556", x"557", x"558",
        x"559", x"55a", x"55b", x"55c", x"55d", x"55e", x"55f", x"560",
        x"561", x"562", x"563", x"564", x"565", x"566", x"567", x"568",
        x"569", x"56a", x"56b", x"56c", x"56d", x"56e", x"56f", x"570",
        x"571", x"572", x"573", x"574", x"575", x"576", x"577", x"578",
        x"579", x"57a", x"57b", x"57c", x"57d", x"57e", x"57f", x"580",
        x"581", x"582", x"583", x"584", x"585", x"586", x"587", x"588",
        x"589", x"58a", x"58b", x"58c", x"58d", x"58e", x"58f", x"590",
        x"591", x"592", x"593", x"594", x"595", x"596", x"597", x"598",
        x"599", x"59a", x"59b", x"59c", x"59d", x"59e", x"59f", x"5a0",
        x"5a1", x"5a2", x"5a3", x"5a4", x"5a5", x"5a6", x"5a7", x"5a8",
        x"5a9", x"5aa", x"5ab", x"5ac", x"5ad", x"5ae", x"5af", x"5b0",
        x"5b1", x"5b2", x"5b3", x"5b4", x"5b5", x"5b6", x"5b7", x"5b8",
        x"5b9", x"5ba", x"5bb", x"5bc", x"5bd", x"5be", x"5bf", x"5c0",
        x"5c1", x"5c2", x"5c3", x"5c4", x"5c5", x"5c6", x"5c7", x"5c8",
        x"5c9", x"5ca", x"5cb", x"5cc", x"5cd", x"5ce", x"5cf", x"5d0",
        x"5d1", x"5d2", x"5d3", x"5d4", x"5d5", x"5d6", x"5d7", x"5d8",
        x"5d9", x"5da", x"5db", x"5dc", x"5dd", x"5de", x"5df", x"5e0",
        x"5e1", x"5e2", x"5e3", x"5e4", x"5e5", x"5e6", x"5e7", x"5e8",
        x"5e9", x"5ea", x"5eb", x"5ec", x"5ed", x"5ee", x"5ef", x"5f0",
        x"5f1", x"5f2", x"5f3", x"5f4", x"5f5", x"5f6", x"5f7", x"5f8",
        x"5f9", x"5fa", x"5fb", x"5fc", x"5fd", x"5fe", x"5ff", x"600",
        x"601", x"602", x"603", x"604", x"605", x"606", x"607", x"608",
        x"609", x"60a", x"60b", x"60c", x"60d", x"60e", x"60f", x"610",
        x"611", x"612", x"613", x"614", x"615", x"616", x"617", x"618",
        x"619", x"61a", x"61b", x"61c", x"61d", x"61e", x"61f", x"620",
        x"621", x"622", x"623", x"624", x"625", x"626", x"627", x"628",
        x"629", x"62a", x"62b", x"62c", x"62d", x"62e", x"62f", x"630",
        x"631", x"632", x"633", x"634", x"635", x"636", x"637", x"638",
        x"639", x"63a", x"63b", x"63c", x"63d", x"63e", x"63f", x"640",
        x"641", x"642", x"643", x"644", x"645", x"646", x"647", x"648",
        x"649", x"64a", x"64b", x"64c", x"64d", x"64e", x"64f", x"650",
        x"651", x"652", x"653", x"654", x"655", x"656", x"657", x"658",
        x"659", x"65a", x"65b", x"65c", x"65d", x"65e", x"65f", x"660",
        x"661", x"662", x"663", x"664", x"665", x"666", x"667", x"668",
        x"669", x"66a", x"66b", x"66c", x"66d", x"66e", x"66f", x"670",
        x"671", x"672", x"673", x"674", x"675", x"676", x"677", x"678",
        x"679", x"67a", x"67b", x"67c", x"67d", x"67e", x"67f", x"680",
        x"681", x"682", x"683", x"684", x"685", x"686", x"687", x"688",
        x"689", x"68a", x"68b", x"68c", x"68d", x"68e", x"68f", x"690",
        x"691", x"692", x"693", x"694", x"695", x"696", x"697", x"698",
        x"699", x"69a", x"69b", x"69c", x"69d", x"69e", x"69f", x"6a0",
        x"6a1", x"6a2", x"6a3", x"6a4", x"6a5", x"6a6", x"6a7", x"6a8",
        x"6a9", x"6aa", x"6ab", x"6ac", x"6ad", x"6ae", x"6af", x"6b0",
        x"6b1", x"6b2", x"6b3", x"6b4", x"6b5", x"6b6", x"6b7", x"6b8",
        x"6b9", x"6ba", x"6bb", x"6bc", x"6bd", x"6be", x"6bf", x"6c0",
        x"6c1", x"6c2", x"6c3", x"6c4", x"6c5", x"6c6", x"6c7", x"6c8",
        x"6c9", x"6ca", x"6cb", x"6cc", x"6cd", x"6ce", x"6cf", x"6d0",
        x"6d1", x"6d2", x"6d3", x"6d4", x"6d5", x"6d6", x"6d7", x"6d8",
        x"6d9", x"6da", x"6db", x"6dc", x"6dd", x"6de", x"6df", x"6e0",
        x"6e1", x"6e2", x"6e3", x"6e4", x"6e5", x"6e6", x"6e7", x"6e8",
        x"6e9", x"6ea", x"6eb", x"6ec", x"6ed", x"6ee", x"6ef", x"6f0",
        x"6f1", x"6f2", x"6f3", x"6f4", x"6f5", x"6f6", x"6f7", x"6f8",
        x"6f9", x"6fa", x"6fb", x"6fc", x"6fd", x"6fe", x"6ff", x"700",
        x"701", x"702", x"703", x"704", x"705", x"706", x"707", x"708",
        x"709", x"70a", x"70b", x"70c", x"70d", x"70e", x"70f", x"710",
        x"711", x"712", x"713", x"714", x"715", x"716", x"717", x"718",
        x"719", x"71a", x"71b", x"71c", x"71d", x"71e", x"71f", x"720",
        x"721", x"722", x"723", x"724", x"725", x"726", x"727", x"728",
        x"729", x"72a", x"72b", x"72c", x"72d", x"72e", x"72f", x"730",
        x"731", x"732", x"733", x"734", x"735", x"736", x"737", x"738",
        x"739", x"73a", x"73b", x"73c", x"73d", x"73e", x"73f", x"740",
        x"741", x"742", x"743", x"744", x"745", x"746", x"747", x"748",
        x"749", x"74a", x"74b", x"74c", x"74d", x"74e", x"74f", x"750",
        x"751", x"752", x"753", x"754", x"755", x"756", x"757", x"758",
        x"759", x"75a", x"75b", x"75c", x"75d", x"75e", x"75f", x"760",
        x"761", x"762", x"763", x"764", x"765", x"766", x"767", x"768",
        x"769", x"76a", x"76b", x"76c", x"76d", x"76e", x"76f", x"770",
        x"771", x"772", x"773", x"774", x"775", x"776", x"777", x"778",
        x"779", x"77a", x"77b", x"77c", x"77d", x"77e", x"77f", x"780",
        x"781", x"782", x"783", x"784", x"785", x"786", x"787", x"788",
        x"789", x"78a", x"78b", x"78c", x"78d", x"78e", x"78f", x"790",
        x"791", x"792", x"793", x"794", x"795", x"796", x"797", x"798",
        x"799", x"79a", x"79b", x"79c", x"79d", x"79e", x"79f", x"7a0",
        x"7a1", x"7a2", x"7a3", x"7a4", x"7a5", x"7a6", x"7a7", x"7a8",
        x"7a9", x"7aa", x"7ab", x"7ac", x"7ad", x"7ae", x"7af", x"7b0",
        x"7b1", x"7b2", x"7b3", x"7b4", x"7b5", x"7b6", x"7b7", x"7b8",
        x"7b9", x"7ba", x"7bb", x"7bc", x"7bd", x"7be", x"7bf", x"7c0",
        x"7c1", x"7c2", x"7c3", x"7c4", x"7c5", x"7c6", x"7c7", x"7c8",
        x"7c9", x"7ca", x"7cb", x"7cc", x"7cd", x"7ce", x"7cf", x"7d0",
        x"7d1", x"7d2", x"7d3", x"7d4", x"7d5", x"7d6", x"7d7", x"7d8",
        x"7d9", x"7da", x"7db", x"7dc", x"7dd", x"7de", x"7df", x"7e0",
        x"7e1", x"7e2", x"7e3", x"7e4", x"7e5", x"7e6", x"7e7", x"7e8",
        x"7e9", x"7ea", x"7eb", x"7ec", x"7ed", x"7ee", x"7ef", x"7f0",
        x"7f1", x"7f2", x"7f3", x"7f4", x"7f5", x"7f6", x"7f7", x"7f8",
        x"7f9", x"7fa", x"7fb", x"7fc", x"7fd", x"7fe", x"7ff", x"800",
        x"801", x"802", x"803", x"804", x"805", x"806", x"807", x"808",
        x"809", x"80a", x"80b", x"80c", x"80d", x"80e", x"80f", x"810",
        x"811", x"812", x"813", x"814", x"815", x"816", x"817", x"818",
        x"819", x"81a", x"81b", x"81c", x"81d", x"81e", x"81f", x"820",
        x"821", x"822", x"823", x"824", x"825", x"826", x"827", x"828",
        x"829", x"82a", x"82b", x"82c", x"82d", x"82e", x"82f", x"830",
        x"831", x"832", x"833", x"834", x"835", x"836", x"837", x"838",
        x"839", x"83a", x"83b", x"83c", x"83d", x"83e", x"83f", x"840",
        x"841", x"842", x"843", x"844", x"845", x"846", x"847", x"848",
        x"849", x"84a", x"84b", x"84c", x"84d", x"84e", x"84f", x"850",
        x"851", x"852", x"853", x"854", x"855", x"856", x"857", x"858",
        x"859", x"85a", x"85b", x"85c", x"85d", x"85e", x"85f", x"860",
        x"861", x"862", x"863", x"864", x"865", x"866", x"867", x"868",
        x"869", x"86a", x"86b", x"86c", x"86d", x"86e", x"86f", x"870",
        x"871", x"872", x"873", x"874", x"875", x"876", x"877", x"878",
        x"879", x"87a", x"87b", x"87c", x"87d", x"87e", x"87f", x"880",
        x"881", x"882", x"883", x"884", x"885", x"886", x"887", x"888",
        x"889", x"88a", x"88b", x"88c", x"88d", x"88e", x"88f", x"890",
        x"891", x"892", x"893", x"894", x"895", x"896", x"897", x"898",
        x"899", x"89a", x"89b", x"89c", x"89d", x"89e", x"89f", x"8a0",
        x"8a1", x"8a2", x"8a3", x"8a4", x"8a5", x"8a6", x"8a7", x"8a8",
        x"8a9", x"8aa", x"8ab", x"8ac", x"8ad", x"8ae", x"8af", x"8b0",
        x"8b1", x"8b2", x"8b3", x"8b4", x"8b5", x"8b6", x"8b7", x"8b8",
        x"8b9", x"8ba", x"8bb", x"8bc", x"8bd", x"8be", x"8bf", x"8c0",
        x"8c1", x"8c2", x"8c3", x"8c4", x"8c5", x"8c6", x"8c7", x"8c8",
        x"8c9", x"8ca", x"8cb", x"8cc", x"8cd", x"8ce", x"8cf", x"8d0",
        x"8d1", x"8d2", x"8d3", x"8d4", x"8d5", x"8d6", x"8d7", x"8d8",
        x"8d9", x"8da", x"8db", x"8dc", x"8dd", x"8de", x"8df", x"8e0",
        x"8e1", x"8e2", x"8e3", x"8e4", x"8e5", x"8e6", x"8e7", x"8e8",
        x"8e9", x"8ea", x"8eb", x"8ec", x"8ed", x"8ee", x"8ef", x"8f0",
        x"8f1", x"8f2", x"8f3", x"8f4", x"8f5", x"8f6", x"8f7", x"8f8",
        x"8f9", x"8fa", x"8fb", x"8fc", x"8fd", x"8fe", x"8ff", x"900",
        x"901", x"902", x"903", x"904", x"905", x"906", x"907", x"908",
        x"909", x"90a", x"90b", x"90c", x"90d", x"90e", x"90f", x"910",
        x"911", x"912", x"913", x"914", x"915", x"916", x"917", x"918",
        x"919", x"91a", x"91b", x"91c", x"91d", x"91e", x"91f", x"920",
        x"921", x"922", x"923", x"924", x"925", x"926", x"927", x"928",
        x"929", x"92a", x"92b", x"92c", x"92d", x"92e", x"92f", x"930",
        x"931", x"932", x"933", x"934", x"935", x"936", x"937", x"938",
        x"939", x"93a", x"93b", x"93c", x"93d", x"93e", x"93f", x"940",
        x"941", x"942", x"943", x"944", x"945", x"946", x"947", x"948",
        x"949", x"94a", x"94b", x"94c", x"94d", x"94e", x"94f", x"950",
        x"951", x"952", x"953", x"954", x"955", x"956", x"957", x"958",
        x"959", x"95a", x"95b", x"95c", x"95d", x"95e", x"95f", x"960",
        x"961", x"962", x"963", x"964", x"965", x"966", x"967", x"968",
        x"969", x"96a", x"96b", x"96c", x"96d", x"96e", x"96f", x"970",
        x"971", x"972", x"973", x"974", x"975", x"976", x"977", x"978",
        x"979", x"97a", x"97b", x"97c", x"97d", x"97e", x"97f", x"980",
        x"981", x"982", x"983", x"984", x"985", x"986", x"987", x"988",
        x"989", x"98a", x"98b", x"98c", x"98d", x"98e", x"98f", x"990",
        x"991", x"992", x"993", x"994", x"995", x"996", x"997", x"998",
        x"999", x"99a", x"99b", x"99c", x"99d", x"99e", x"99f", x"9a0",
        x"9a1", x"9a2", x"9a3", x"9a4", x"9a5", x"9a6", x"9a7", x"9a8",
        x"9a9", x"9aa", x"9ab", x"9ac", x"9ad", x"9ae", x"9af", x"9b0",
        x"9b1", x"9b2", x"9b3", x"9b4", x"9b5", x"9b6", x"9b7", x"9b8",
        x"9b9", x"9ba", x"9bb", x"9bc", x"9bd", x"9be", x"9bf", x"9c0",
        x"9c1", x"9c2", x"9c3", x"9c4", x"9c5", x"9c6", x"9c7", x"9c8",
        x"9c9", x"9ca", x"9cb", x"9cc", x"9cd", x"9ce", x"9cf", x"9d0",
        x"9d1", x"9d2", x"9d3", x"9d4", x"9d5", x"9d6", x"9d7", x"9d8",
        x"9d9", x"9da", x"9db", x"9dc", x"9dd", x"9de", x"9df", x"9e0",
        x"9e1", x"9e2", x"9e3", x"9e4", x"9e5", x"9e6", x"9e7", x"9e8",
        x"9e9", x"9ea", x"9eb", x"9ec", x"9ed", x"9ee", x"9ef", x"9f0",
        x"9f1", x"9f2", x"9f3", x"9f4", x"9f5", x"9f6", x"9f7", x"9f8",
        x"9f9", x"9fa", x"9fb", x"9fc", x"9fd", x"9fe", x"9ff", x"a00",
        x"a01", x"a02", x"a03", x"a04", x"a05", x"a06", x"a07", x"a08",
        x"a09", x"a0a", x"a0b", x"a0c", x"a0d", x"a0e", x"a0f", x"a10",
        x"a11", x"a12", x"a13", x"a14", x"a15", x"a16", x"a17", x"a18",
        x"a19", x"a1a", x"a1b", x"a1c", x"a1d", x"a1e", x"a1f", x"a20",
        x"a21", x"a22", x"a23", x"a24", x"a25", x"a26", x"a27", x"a28",
        x"a29", x"a2a", x"a2b", x"a2c", x"a2d", x"a2e", x"a2f", x"a30",
        x"a31", x"a32", x"a33", x"a34", x"a35", x"a36", x"a37", x"a38",
        x"a39", x"a3a", x"a3b", x"a3c", x"a3d", x"a3e", x"a3f", x"a40",
        x"a41", x"a42", x"a43", x"a44", x"a45", x"a46", x"a47", x"a48",
        x"a49", x"a4a", x"a4b", x"a4c", x"a4d", x"a4e", x"a4f", x"a50",
        x"a51", x"a52", x"a53", x"a54", x"a55", x"a56", x"a57", x"a58",
        x"a59", x"a5a", x"a5b", x"a5c", x"a5d", x"a5e", x"a5f", x"a60",
        x"a61", x"a62", x"a63", x"a64", x"a65", x"a66", x"a67", x"a68",
        x"a69", x"a6a", x"a6b", x"a6c", x"a6d", x"a6e", x"a6f", x"a70",
        x"a71", x"a72", x"a73", x"a74", x"a75", x"a76", x"a77", x"a78",
        x"a79", x"a7a", x"a7b", x"a7c", x"a7d", x"a7e", x"a7f", x"a80",
        x"a81", x"a82", x"a83", x"a84", x"a85", x"a86", x"a87", x"a88",
        x"a89", x"a8a", x"a8b", x"a8c", x"a8d", x"a8e", x"a8f", x"a90",
        x"a91", x"a92", x"a93", x"a94", x"a95", x"a96", x"a97", x"a98",
        x"a99", x"a9a", x"a9b", x"a9c", x"a9d", x"a9e", x"a9f", x"aa0",
        x"aa1", x"aa2", x"aa3", x"aa4", x"aa5", x"aa6", x"aa7", x"aa8",
        x"aa9", x"aaa", x"aab", x"aac", x"aad", x"aae", x"aaf", x"ab0",
        x"ab1", x"ab2", x"ab3", x"ab4", x"ab5", x"ab6", x"ab7", x"ab8",
        x"ab9", x"aba", x"abb", x"abc", x"abd", x"abe", x"abf", x"ac0",
        x"ac1", x"ac2", x"ac3", x"ac4", x"ac5", x"ac6", x"ac7", x"ac8",
        x"ac9", x"aca", x"acb", x"acc", x"acd", x"ace", x"acf", x"ad0",
        x"ad1", x"ad2", x"ad3", x"ad4", x"ad5", x"ad6", x"ad7", x"ad8",
        x"ad9", x"ada", x"adb", x"adc", x"add", x"ade", x"adf", x"ae0",
        x"ae1", x"ae2", x"ae3", x"ae4", x"ae5", x"ae6", x"ae7", x"ae8",
        x"ae9", x"aea", x"aeb", x"aec", x"aed", x"aee", x"aef", x"af0",
        x"af1", x"af2", x"af3", x"af4", x"af5", x"af6", x"af7", x"af8",
        x"af9", x"afa", x"afb", x"afc", x"afd", x"afe", x"aff", x"b00",
        x"b01", x"b02", x"b03", x"b04", x"b05", x"b06", x"b07", x"b08",
        x"b09", x"b0a", x"b0b", x"b0c", x"b0d", x"b0e", x"b0f", x"b10",
        x"b11", x"b12", x"b13", x"b14", x"b15", x"b16", x"b17", x"b18",
        x"b19", x"b1a", x"b1b", x"b1c", x"b1d", x"b1e", x"b1f", x"b20",
        x"b21", x"b22", x"b23", x"b24", x"b25", x"b26", x"b27", x"b28",
        x"b29", x"b2a", x"b2b", x"b2c", x"b2d", x"b2e", x"b2f", x"b30",
        x"b31", x"b32", x"b33", x"b34", x"b35", x"b36", x"b37", x"b38",
        x"b39", x"b3a", x"b3b", x"b3c", x"b3d", x"b3e", x"b3f", x"b40",
        x"b41", x"b42", x"b43", x"b44", x"b45", x"b46", x"b47", x"b48",
        x"b49", x"b4a", x"b4b", x"b4c", x"b4d", x"b4e", x"b4f", x"b50",
        x"b51", x"b52", x"b53", x"b54", x"b55", x"b56", x"b57", x"b58",
        x"b59", x"b5a", x"b5b", x"b5c", x"b5d", x"b5e", x"b5f", x"b60",
        x"b61", x"b62", x"b63", x"b64", x"b65", x"b66", x"b67", x"b68",
        x"b69", x"b6a", x"b6b", x"b6c", x"b6d", x"b6e", x"b6f", x"b70",
        x"b71", x"b72", x"b73", x"b74", x"b75", x"b76", x"b77", x"b78",
        x"b79", x"b7a", x"b7b", x"b7c", x"b7d", x"b7e", x"b7f", x"b80",
        x"b81", x"b82", x"b83", x"b84", x"b85", x"b86", x"b87", x"b88",
        x"b89", x"b8a", x"b8b", x"b8c", x"b8d", x"b8e", x"b8f", x"b90",
        x"b91", x"b92", x"b93", x"b94", x"b95", x"b96", x"b97", x"b98",
        x"b99", x"b9a", x"b9b", x"b9c", x"b9d", x"b9e", x"b9f", x"ba0",
        x"ba1", x"ba2", x"ba3", x"ba4", x"ba5", x"ba6", x"ba7", x"ba8",
        x"ba9", x"baa", x"bab", x"bac", x"bad", x"bae", x"baf", x"bb0",
        x"bb1", x"bb2", x"bb3", x"bb4", x"bb5", x"bb6", x"bb7", x"bb8",
        x"bb9", x"bba", x"bbb", x"bbc", x"bbd", x"bbe", x"bbf", x"bc0",
        x"bc1", x"bc2", x"bc3", x"bc4", x"bc5", x"bc6", x"bc7", x"bc8",
        x"bc9", x"bca", x"bcb", x"bcc", x"bcd", x"bce", x"bcf", x"bd0",
        x"bd1", x"bd2", x"bd3", x"bd4", x"bd5", x"bd6", x"bd7", x"bd8",
        x"bd9", x"bda", x"bdb", x"bdc", x"bdd", x"bde", x"bdf", x"be0",
        x"be1", x"be2", x"be3", x"be4", x"be5", x"be6", x"be7", x"be8",
        x"be9", x"bea", x"beb", x"bec", x"bed", x"bee", x"bef", x"bf0",
        x"bf1", x"bf2", x"bf3", x"bf4", x"bf5", x"bf6", x"bf7", x"bf8",
        x"bf9", x"bfa", x"bfb", x"bfc", x"bfd", x"bfe", x"bff", x"c00",
        x"c01", x"c02", x"c03", x"c04", x"c05", x"c06", x"c07", x"c08",
        x"c09", x"c0a", x"c0b", x"c0c", x"c0d", x"c0e", x"c0f", x"c10",
        x"c11", x"c12", x"c13", x"c14", x"c15", x"c16", x"c17", x"c18",
        x"c19", x"c1a", x"c1b", x"c1c", x"c1d", x"c1e", x"c1f", x"c20",
        x"c21", x"c22", x"c23", x"c24", x"c25", x"c26", x"c27", x"c28",
        x"c29", x"c2a", x"c2b", x"c2c", x"c2d", x"c2e", x"c2f", x"c30",
        x"c31", x"c32", x"c33", x"c34", x"c35", x"c36", x"c37", x"c38",
        x"c39", x"c3a", x"c3b", x"c3c", x"c3d", x"c3e", x"c3f", x"c40",
        x"c41", x"c42", x"c43", x"c44", x"c45", x"c46", x"c47", x"c48",
        x"c49", x"c4a", x"c4b", x"c4c", x"c4d", x"c4e", x"c4f", x"c50",
        x"c51", x"c52", x"c53", x"c54", x"c55", x"c56", x"c57", x"c58",
        x"c59", x"c5a", x"c5b", x"c5c", x"c5d", x"c5e", x"c5f", x"c60",
        x"c61", x"c62", x"c63", x"c64", x"c65", x"c66", x"c67", x"c68",
        x"c69", x"c6a", x"c6b", x"c6c", x"c6d", x"c6e", x"c6f", x"c70",
        x"c71", x"c72", x"c73", x"c74", x"c75", x"c76", x"c77", x"c78",
        x"c79", x"c7a", x"c7b", x"c7c", x"c7d", x"c7e", x"c7f", x"c80",
        x"c81", x"c82", x"c83", x"c84", x"c85", x"c86", x"c87", x"c88",
        x"c89", x"c8a", x"c8b", x"c8c", x"c8d", x"c8e", x"c8f", x"c90",
        x"c91", x"c92", x"c93", x"c94", x"c95", x"c96", x"c97", x"c98",
        x"c99", x"c9a", x"c9b", x"c9c", x"c9d", x"c9e", x"c9f", x"ca0",
        x"ca1", x"ca2", x"ca3", x"ca4", x"ca5", x"ca6", x"ca7", x"ca8",
        x"ca9", x"caa", x"cab", x"cac", x"cad", x"cae", x"caf", x"cb0",
        x"cb1", x"cb2", x"cb3", x"cb4", x"cb5", x"cb6", x"cb7", x"cb8",
        x"cb9", x"cba", x"cbb", x"cbc", x"cbd", x"cbe", x"cbf", x"cc0",
        x"cc1", x"cc2", x"cc3", x"cc4", x"cc5", x"cc6", x"cc7", x"cc8",
        x"cc9", x"cca", x"ccb", x"ccc", x"ccd", x"cce", x"ccf", x"cd0",
        x"cd1", x"cd2", x"cd3", x"cd4", x"cd5", x"cd6", x"cd7", x"cd8",
        x"cd9", x"cda", x"cdb", x"cdc", x"cdd", x"cde", x"cdf", x"ce0",
        x"ce1", x"ce2", x"ce3", x"ce4", x"ce5", x"ce6", x"ce7", x"ce8",
        x"ce9", x"cea", x"ceb", x"cec", x"ced", x"cee", x"cef", x"cf0",
        x"cf1", x"cf2", x"cf3", x"cf4", x"cf5", x"cf6", x"cf7", x"cf8",
        x"cf9", x"cfa", x"cfb", x"cfc", x"cfd", x"cfe", x"cff", x"d00",
        x"d01", x"d02", x"d03", x"d04", x"d05", x"d06", x"d07", x"d08",
        x"d09", x"d0a", x"d0b", x"d0c", x"d0d", x"d0e", x"d0f", x"d10",
        x"d11", x"d12", x"d13", x"d14", x"d15", x"d16", x"d17", x"d18",
        x"d19", x"d1a", x"d1b", x"d1c", x"d1d", x"d1e", x"d1f", x"d20",
        x"d21", x"d22", x"d23", x"d24", x"d25", x"d26", x"d27", x"d28",
        x"d29", x"d2a", x"d2b", x"d2c", x"d2d", x"d2e", x"d2f", x"d30",
        x"d31", x"d32", x"d33", x"d34", x"d35", x"d36", x"d37", x"d38",
        x"d39", x"d3a", x"d3b", x"d3c", x"d3d", x"d3e", x"d3f", x"d40",
        x"d41", x"d42", x"d43", x"d44", x"d45", x"d46", x"d47", x"d48",
        x"d49", x"d4a", x"d4b", x"d4c", x"d4d", x"d4e", x"d4f", x"d50",
        x"d51", x"d52", x"d53", x"d54", x"d55", x"d56", x"d57", x"d58",
        x"d59", x"d5a", x"d5b", x"d5c", x"d5d", x"d5e", x"d5f", x"d60",
        x"d61", x"d62", x"d63", x"d64", x"d65", x"d66", x"d67", x"d68",
        x"d69", x"d6a", x"d6b", x"d6c", x"d6d", x"d6e", x"d6f", x"d70",
        x"d71", x"d72", x"d73", x"d74", x"d75", x"d76", x"d77", x"d78",
        x"d79", x"d7a", x"d7b", x"d7c", x"d7d", x"d7e", x"d7f", x"d80",
        x"d81", x"d82", x"d83", x"d84", x"d85", x"d86", x"d87", x"d88",
        x"d89", x"d8a", x"d8b", x"d8c", x"d8d", x"d8e", x"d8f", x"d90",
        x"d91", x"d92", x"d93", x"d94", x"d95", x"d96", x"d97", x"d98",
        x"d99", x"d9a", x"d9b", x"d9c", x"d9d", x"d9e", x"d9f", x"da0",
        x"da1", x"da2", x"da3", x"da4", x"da5", x"da6", x"da7", x"da8",
        x"da9", x"daa", x"dab", x"dac", x"dad", x"dae", x"daf", x"db0",
        x"db1", x"db2", x"db3", x"db4", x"db5", x"db6", x"db7", x"db8",
        x"db9", x"dba", x"dbb", x"dbc", x"dbd", x"dbe", x"dbf", x"dc0",
        x"dc1", x"dc2", x"dc3", x"dc4", x"dc5", x"dc6", x"dc7", x"dc8",
        x"dc9", x"dca", x"dcb", x"dcc", x"dcd", x"dce", x"dcf", x"dd0",
        x"dd1", x"dd2", x"dd3", x"dd4", x"dd5", x"dd6", x"dd7", x"dd8",
        x"dd9", x"dda", x"ddb", x"ddc", x"ddd", x"dde", x"ddf", x"de0",
        x"de1", x"de2", x"de3", x"de4", x"de5", x"de6", x"de7", x"de8",
        x"de9", x"dea", x"deb", x"dec", x"ded", x"dee", x"def", x"df0",
        x"df1", x"df2", x"df3", x"df4", x"df5", x"df6", x"df7", x"df8",
        x"df9", x"dfa", x"dfb", x"dfc", x"dfd", x"dfe", x"dff", x"e00",
        x"e01", x"e02", x"e03", x"e04", x"e05", x"e06", x"e07", x"e08",
        x"e09", x"e0a", x"e0b", x"e0c", x"e0d", x"e0e", x"e0f", x"e10",
        x"e11", x"e12", x"e13", x"e14", x"e15", x"e16", x"e17", x"e18",
        x"e19", x"e1a", x"e1b", x"e1c", x"e1d", x"e1e", x"e1f", x"e20",
        x"e21", x"e22", x"e23", x"e24", x"e25", x"e26", x"e27", x"e28",
        x"e29", x"e2a", x"e2b", x"e2c", x"e2d", x"e2e", x"e2f", x"e30",
        x"e31", x"e32", x"e33", x"e34", x"e35", x"e36", x"e37", x"e38",
        x"e39", x"e3a", x"e3b", x"e3c", x"e3d", x"e3e", x"e3f", x"e40",
        x"e41", x"e42", x"e43", x"e44", x"e45", x"e46", x"e47", x"e48",
        x"e49", x"e4a", x"e4b", x"e4c", x"e4d", x"e4e", x"e4f", x"e50",
        x"e51", x"e52", x"e53", x"e54", x"e55", x"e56", x"e57", x"e58",
        x"e59", x"e5a", x"e5b", x"e5c", x"e5d", x"e5e", x"e5f", x"e60",
        x"e61", x"e62", x"e63", x"e64", x"e65", x"e66", x"e67", x"e68",
        x"e69", x"e6a", x"e6b", x"e6c", x"e6d", x"e6e", x"e6f", x"e70",
        x"e71", x"e72", x"e73", x"e74", x"e75", x"e76", x"e77", x"e78",
        x"e79", x"e7a", x"e7b", x"e7c", x"e7d", x"e7e", x"e7f", x"e80",
        x"e81", x"e82", x"e83", x"e84", x"e85", x"e86", x"e87", x"e88",
        x"e89", x"e8a", x"e8b", x"e8c", x"e8d", x"e8e", x"e8f", x"e90",
        x"e91", x"e92", x"e93", x"e94", x"e95", x"e96", x"e97", x"e98",
        x"e99", x"e9a", x"e9b", x"e9c", x"e9d", x"e9e", x"e9f", x"ea0",
        x"ea1", x"ea2", x"ea3", x"ea4", x"ea5", x"ea6", x"ea7", x"ea8",
        x"ea9", x"eaa", x"eab", x"eac", x"ead", x"eae", x"eaf", x"eb0",
        x"eb1", x"eb2", x"eb3", x"eb4", x"eb5", x"eb6", x"eb7", x"eb8",
        x"eb9", x"eba", x"ebb", x"ebc", x"ebd", x"ebe", x"ebf", x"ec0",
        x"ec1", x"ec2", x"ec3", x"ec4", x"ec5", x"ec6", x"ec7", x"ec8",
        x"ec9", x"eca", x"ecb", x"ecc", x"ecd", x"ece", x"ecf", x"ed0",
        x"ed1", x"ed2", x"ed3", x"ed4", x"ed5", x"ed6", x"ed7", x"ed8",
        x"ed9", x"eda", x"edb", x"edc", x"edd", x"ede", x"edf", x"ee0",
        x"ee1", x"ee2", x"ee3", x"ee4", x"ee5", x"ee6", x"ee7", x"ee8",
        x"ee9", x"eea", x"eeb", x"eec", x"eed", x"eee", x"eef", x"ef0",
        x"ef1", x"ef2", x"ef3", x"ef4", x"ef5", x"ef6", x"ef7", x"ef8",
        x"ef9", x"efa", x"efb", x"efc", x"efd", x"efe", x"eff", x"f00",
        x"f01", x"f02", x"f03", x"f04", x"f05", x"f06", x"f07", x"f08",
        x"f09", x"f0a", x"f0b", x"f0c", x"f0d", x"f0e", x"f0f", x"f10",
        x"f11", x"f12", x"f13", x"f14", x"f15", x"f16", x"f17", x"f18",
        x"f19", x"f1a", x"f1b", x"f1c", x"f1d", x"f1e", x"f1f", x"f20",
        x"f21", x"f22", x"f23", x"f24", x"f25", x"f26", x"f27", x"f28",
        x"f29", x"f2a", x"f2b", x"f2c", x"f2d", x"f2e", x"f2f", x"f30",
        x"f31", x"f32", x"f33", x"f34", x"f35", x"f36", x"f37", x"f38",
        x"f39", x"f3a", x"f3b", x"f3c", x"f3d", x"f3e", x"f3f", x"f40",
        x"f41", x"f42", x"f43", x"f44", x"f45", x"f46", x"f47", x"f48",
        x"f49", x"f4a", x"f4b", x"f4c", x"f4d", x"f4e", x"f4f", x"f50",
        x"f51", x"f52", x"f53", x"f54", x"f55", x"f56", x"f57", x"f58",
        x"f59", x"f5a", x"f5b", x"f5c", x"f5d", x"f5e", x"f5f", x"f60",
        x"f61", x"f62", x"f63", x"f64", x"f65", x"f66", x"f67", x"f68",
        x"f69", x"f6a", x"f6b", x"f6c", x"f6d", x"f6e", x"f6f", x"f70",
        x"f71", x"f72", x"f73", x"f74", x"f75", x"f76", x"f77", x"f78",
        x"f79", x"f7a", x"f7b", x"f7c", x"f7d", x"f7e", x"f7f", x"f80",
        x"f81", x"f82", x"f83", x"f84", x"f85", x"f86", x"f87", x"f88",
        x"f89", x"f8a", x"f8b", x"f8c", x"f8d", x"f8e", x"f8f", x"f90",
        x"f91", x"f92", x"f93", x"f94", x"f95", x"f96", x"f97", x"f98",
        x"f99", x"f9a", x"f9b", x"f9c", x"f9d", x"f9e", x"f9f", x"fa0",
        x"fa1", x"fa2", x"fa3", x"fa4", x"fa5", x"fa6", x"fa7", x"fa8",
        x"fa9", x"faa", x"fab", x"fac", x"fad", x"fae", x"faf", x"fb0",
        x"fb1", x"fb2", x"fb3", x"fb4", x"fb5", x"fb6", x"fb7", x"fb8",
        x"fb9", x"fba", x"fbb", x"fbc", x"fbd", x"fbe", x"fbf", x"fc0",
        x"fc1", x"fc2", x"fc3", x"fc4", x"fc5", x"fc6", x"fc7", x"fc8",
        x"fc9", x"fca", x"fcb", x"fcc", x"fcd", x"fce", x"fcf", x"fd0",
        x"fd1", x"fd2", x"fd3", x"fd4", x"fd5", x"fd6", x"fd7", x"fd8",
        x"fd9", x"fda", x"fdb", x"fdc", x"fdd", x"fde", x"fdf", x"fe0",
        x"fe1", x"fe2", x"fe3", x"fe4", x"fe5", x"fe6", x"fe7", x"fe8",
        x"fe9", x"fea", x"feb", x"fec", x"fed", x"fee", x"fef", x"ff0",
        x"ff1", x"ff2", x"ff3", x"ff4", x"ff5", x"ff6", x"ff7", x"ff8",
        x"ff9", x"ffa", x"ffb", x"ffc", x"ffd", x"ffe", x"fff", x"000"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr,clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp,en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
