library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(11 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom;

architecture arch of rom is
    type memoria_rom is array (0 to 4095) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"800", x"803", x"806", x"809", x"80c", x"80f", x"812", x"815",
        x"819", x"81c", x"81f", x"822", x"825", x"828", x"82b", x"82f",
        x"832", x"835", x"838", x"83b", x"83e", x"841", x"845", x"848",
        x"84b", x"84e", x"851", x"854", x"857", x"85b", x"85e", x"861",
        x"864", x"867", x"86a", x"86d", x"871", x"874", x"877", x"87a",
        x"87d", x"880", x"883", x"886", x"88a", x"88d", x"890", x"893",
        x"896", x"899", x"89c", x"8a0", x"8a3", x"8a6", x"8a9", x"8ac",
        x"8af", x"8b2", x"8b5", x"8b9", x"8bc", x"8bf", x"8c2", x"8c5",
        x"8c8", x"8cb", x"8ce", x"8d2", x"8d5", x"8d8", x"8db", x"8de",
        x"8e1", x"8e4", x"8e7", x"8eb", x"8ee", x"8f1", x"8f4", x"8f7",
        x"8fa", x"8fd", x"900", x"903", x"907", x"90a", x"90d", x"910",
        x"913", x"916", x"919", x"91c", x"91f", x"923", x"926", x"929",
        x"92c", x"92f", x"932", x"935", x"938", x"93b", x"93f", x"942",
        x"945", x"948", x"94b", x"94e", x"951", x"954", x"957", x"95a",
        x"95e", x"961", x"964", x"967", x"96a", x"96d", x"970", x"973",
        x"976", x"979", x"97c", x"980", x"983", x"986", x"989", x"98c",
        x"98f", x"992", x"995", x"998", x"99b", x"99e", x"9a1", x"9a4",
        x"9a8", x"9ab", x"9ae", x"9b1", x"9b4", x"9b7", x"9ba", x"9bd",
        x"9c0", x"9c3", x"9c6", x"9c9", x"9cc", x"9cf", x"9d2", x"9d6",
        x"9d9", x"9dc", x"9df", x"9e2", x"9e5", x"9e8", x"9eb", x"9ee",
        x"9f1", x"9f4", x"9f7", x"9fa", x"9fd", x"a00", x"a03", x"a06",
        x"a09", x"a0c", x"a0f", x"a12", x"a15", x"a19", x"a1c", x"a1f",
        x"a22", x"a25", x"a28", x"a2b", x"a2e", x"a31", x"a34", x"a37",
        x"a3a", x"a3d", x"a40", x"a43", x"a46", x"a49", x"a4c", x"a4f",
        x"a52", x"a55", x"a58", x"a5b", x"a5e", x"a61", x"a64", x"a67",
        x"a6a", x"a6d", x"a70", x"a73", x"a76", x"a79", x"a7c", x"a7f",
        x"a82", x"a85", x"a88", x"a8b", x"a8e", x"a91", x"a94", x"a97",
        x"a9a", x"a9d", x"aa0", x"aa2", x"aa5", x"aa8", x"aab", x"aae",
        x"ab1", x"ab4", x"ab7", x"aba", x"abd", x"ac0", x"ac3", x"ac6",
        x"ac9", x"acc", x"acf", x"ad2", x"ad5", x"ad8", x"adb", x"add",
        x"ae0", x"ae3", x"ae6", x"ae9", x"aec", x"aef", x"af2", x"af5",
        x"af8", x"afb", x"afe", x"b01", x"b03", x"b06", x"b09", x"b0c",
        x"b0f", x"b12", x"b15", x"b18", x"b1b", x"b1e", x"b20", x"b23",
        x"b26", x"b29", x"b2c", x"b2f", x"b32", x"b35", x"b37", x"b3a",
        x"b3d", x"b40", x"b43", x"b46", x"b49", x"b4c", x"b4e", x"b51",
        x"b54", x"b57", x"b5a", x"b5d", x"b60", x"b62", x"b65", x"b68",
        x"b6b", x"b6e", x"b71", x"b73", x"b76", x"b79", x"b7c", x"b7f",
        x"b82", x"b84", x"b87", x"b8a", x"b8d", x"b90", x"b92", x"b95",
        x"b98", x"b9b", x"b9e", x"ba0", x"ba3", x"ba6", x"ba9", x"bac",
        x"bae", x"bb1", x"bb4", x"bb7", x"bba", x"bbc", x"bbf", x"bc2",
        x"bc5", x"bc7", x"bca", x"bcd", x"bd0", x"bd3", x"bd5", x"bd8",
        x"bdb", x"bde", x"be0", x"be3", x"be6", x"be9", x"beb", x"bee",
        x"bf1", x"bf3", x"bf6", x"bf9", x"bfc", x"bfe", x"c01", x"c04",
        x"c06", x"c09", x"c0c", x"c0f", x"c11", x"c14", x"c17", x"c19",
        x"c1c", x"c1f", x"c22", x"c24", x"c27", x"c2a", x"c2c", x"c2f",
        x"c32", x"c34", x"c37", x"c3a", x"c3c", x"c3f", x"c42", x"c44",
        x"c47", x"c4a", x"c4c", x"c4f", x"c52", x"c54", x"c57", x"c59",
        x"c5c", x"c5f", x"c61", x"c64", x"c67", x"c69", x"c6c", x"c6e",
        x"c71", x"c74", x"c76", x"c79", x"c7b", x"c7e", x"c81", x"c83",
        x"c86", x"c88", x"c8b", x"c8e", x"c90", x"c93", x"c95", x"c98",
        x"c9a", x"c9d", x"ca0", x"ca2", x"ca5", x"ca7", x"caa", x"cac",
        x"caf", x"cb1", x"cb4", x"cb7", x"cb9", x"cbc", x"cbe", x"cc1",
        x"cc3", x"cc6", x"cc8", x"ccb", x"ccd", x"cd0", x"cd2", x"cd5",
        x"cd7", x"cda", x"cdc", x"cdf", x"ce1", x"ce4", x"ce6", x"ce9",
        x"ceb", x"cee", x"cf0", x"cf3", x"cf5", x"cf8", x"cfa", x"cfc",
        x"cff", x"d01", x"d04", x"d06", x"d09", x"d0b", x"d0e", x"d10",
        x"d12", x"d15", x"d17", x"d1a", x"d1c", x"d1f", x"d21", x"d23",
        x"d26", x"d28", x"d2b", x"d2d", x"d2f", x"d32", x"d34", x"d36",
        x"d39", x"d3b", x"d3e", x"d40", x"d42", x"d45", x"d47", x"d49",
        x"d4c", x"d4e", x"d50", x"d53", x"d55", x"d58", x"d5a", x"d5c",
        x"d5f", x"d61", x"d63", x"d65", x"d68", x"d6a", x"d6c", x"d6f",
        x"d71", x"d73", x"d76", x"d78", x"d7a", x"d7c", x"d7f", x"d81",
        x"d83", x"d86", x"d88", x"d8a", x"d8c", x"d8f", x"d91", x"d93",
        x"d95", x"d98", x"d9a", x"d9c", x"d9e", x"da1", x"da3", x"da5",
        x"da7", x"daa", x"dac", x"dae", x"db0", x"db2", x"db5", x"db7",
        x"db9", x"dbb", x"dbd", x"dc0", x"dc2", x"dc4", x"dc6", x"dc8",
        x"dca", x"dcd", x"dcf", x"dd1", x"dd3", x"dd5", x"dd7", x"dd9",
        x"ddc", x"dde", x"de0", x"de2", x"de4", x"de6", x"de8", x"dea",
        x"ded", x"def", x"df1", x"df3", x"df5", x"df7", x"df9", x"dfb",
        x"dfd", x"dff", x"e02", x"e04", x"e06", x"e08", x"e0a", x"e0c",
        x"e0e", x"e10", x"e12", x"e14", x"e16", x"e18", x"e1a", x"e1c",
        x"e1e", x"e20", x"e22", x"e24", x"e26", x"e28", x"e2a", x"e2c",
        x"e2e", x"e30", x"e32", x"e34", x"e36", x"e38", x"e3a", x"e3c",
        x"e3e", x"e40", x"e42", x"e44", x"e46", x"e48", x"e4a", x"e4c",
        x"e4e", x"e50", x"e51", x"e53", x"e55", x"e57", x"e59", x"e5b",
        x"e5d", x"e5f", x"e61", x"e63", x"e65", x"e66", x"e68", x"e6a",
        x"e6c", x"e6e", x"e70", x"e72", x"e74", x"e75", x"e77", x"e79",
        x"e7b", x"e7d", x"e7f", x"e80", x"e82", x"e84", x"e86", x"e88",
        x"e8a", x"e8b", x"e8d", x"e8f", x"e91", x"e92", x"e94", x"e96",
        x"e98", x"e9a", x"e9b", x"e9d", x"e9f", x"ea1", x"ea2", x"ea4",
        x"ea6", x"ea8", x"ea9", x"eab", x"ead", x"eaf", x"eb0", x"eb2",
        x"eb4", x"eb5", x"eb7", x"eb9", x"ebb", x"ebc", x"ebe", x"ec0",
        x"ec1", x"ec3", x"ec5", x"ec6", x"ec8", x"eca", x"ecb", x"ecd",
        x"ecf", x"ed0", x"ed2", x"ed4", x"ed5", x"ed7", x"ed8", x"eda",
        x"edc", x"edd", x"edf", x"ee1", x"ee2", x"ee4", x"ee5", x"ee7",
        x"ee8", x"eea", x"eec", x"eed", x"eef", x"ef0", x"ef2", x"ef3",
        x"ef5", x"ef7", x"ef8", x"efa", x"efb", x"efd", x"efe", x"f00",
        x"f01", x"f03", x"f04", x"f06", x"f07", x"f09", x"f0a", x"f0c",
        x"f0d", x"f0f", x"f10", x"f12", x"f13", x"f15", x"f16", x"f17",
        x"f19", x"f1a", x"f1c", x"f1d", x"f1f", x"f20", x"f22", x"f23",
        x"f24", x"f26", x"f27", x"f29", x"f2a", x"f2b", x"f2d", x"f2e",
        x"f30", x"f31", x"f32", x"f34", x"f35", x"f36", x"f38", x"f39",
        x"f3a", x"f3c", x"f3d", x"f3e", x"f40", x"f41", x"f42", x"f44",
        x"f45", x"f46", x"f48", x"f49", x"f4a", x"f4c", x"f4d", x"f4e",
        x"f4f", x"f51", x"f52", x"f53", x"f54", x"f56", x"f57", x"f58",
        x"f59", x"f5b", x"f5c", x"f5d", x"f5e", x"f60", x"f61", x"f62",
        x"f63", x"f64", x"f66", x"f67", x"f68", x"f69", x"f6a", x"f6b",
        x"f6d", x"f6e", x"f6f", x"f70", x"f71", x"f72", x"f74", x"f75",
        x"f76", x"f77", x"f78", x"f79", x"f7a", x"f7b", x"f7d", x"f7e",
        x"f7f", x"f80", x"f81", x"f82", x"f83", x"f84", x"f85", x"f86",
        x"f87", x"f88", x"f89", x"f8a", x"f8c", x"f8d", x"f8e", x"f8f",
        x"f90", x"f91", x"f92", x"f93", x"f94", x"f95", x"f96", x"f97",
        x"f98", x"f99", x"f9a", x"f9b", x"f9c", x"f9d", x"f9d", x"f9e",
        x"f9f", x"fa0", x"fa1", x"fa2", x"fa3", x"fa4", x"fa5", x"fa6",
        x"fa7", x"fa8", x"fa9", x"faa", x"faa", x"fab", x"fac", x"fad",
        x"fae", x"faf", x"fb0", x"fb1", x"fb1", x"fb2", x"fb3", x"fb4",
        x"fb5", x"fb6", x"fb6", x"fb7", x"fb8", x"fb9", x"fba", x"fbb",
        x"fbb", x"fbc", x"fbd", x"fbe", x"fbf", x"fbf", x"fc0", x"fc1",
        x"fc2", x"fc2", x"fc3", x"fc4", x"fc5", x"fc5", x"fc6", x"fc7",
        x"fc8", x"fc8", x"fc9", x"fca", x"fca", x"fcb", x"fcc", x"fcd",
        x"fcd", x"fce", x"fcf", x"fcf", x"fd0", x"fd1", x"fd1", x"fd2",
        x"fd3", x"fd3", x"fd4", x"fd5", x"fd5", x"fd6", x"fd6", x"fd7",
        x"fd8", x"fd8", x"fd9", x"fd9", x"fda", x"fdb", x"fdb", x"fdc",
        x"fdc", x"fdd", x"fde", x"fde", x"fdf", x"fdf", x"fe0", x"fe0",
        x"fe1", x"fe1", x"fe2", x"fe2", x"fe3", x"fe3", x"fe4", x"fe4",
        x"fe5", x"fe5", x"fe6", x"fe6", x"fe7", x"fe7", x"fe8", x"fe8",
        x"fe9", x"fe9", x"fea", x"fea", x"feb", x"feb", x"fec", x"fec",
        x"fec", x"fed", x"fed", x"fee", x"fee", x"fee", x"fef", x"fef",
        x"ff0", x"ff0", x"ff0", x"ff1", x"ff1", x"ff1", x"ff2", x"ff2",
        x"ff3", x"ff3", x"ff3", x"ff4", x"ff4", x"ff4", x"ff5", x"ff5",
        x"ff5", x"ff5", x"ff6", x"ff6", x"ff6", x"ff7", x"ff7", x"ff7",
        x"ff7", x"ff8", x"ff8", x"ff8", x"ff8", x"ff9", x"ff9", x"ff9",
        x"ff9", x"ffa", x"ffa", x"ffa", x"ffa", x"ffb", x"ffb", x"ffb",
        x"ffb", x"ffb", x"ffc", x"ffc", x"ffc", x"ffc", x"ffc", x"ffc",
        x"ffd", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd",
        x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe",
        x"ffe", x"ffe", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ffe",
        x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe", x"ffe",
        x"ffe", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd", x"ffd",
        x"ffd", x"ffc", x"ffc", x"ffc", x"ffc", x"ffc", x"ffc", x"ffb",
        x"ffb", x"ffb", x"ffb", x"ffb", x"ffa", x"ffa", x"ffa", x"ffa",
        x"ff9", x"ff9", x"ff9", x"ff9", x"ff8", x"ff8", x"ff8", x"ff8",
        x"ff7", x"ff7", x"ff7", x"ff7", x"ff6", x"ff6", x"ff6", x"ff5",
        x"ff5", x"ff5", x"ff5", x"ff4", x"ff4", x"ff4", x"ff3", x"ff3",
        x"ff3", x"ff2", x"ff2", x"ff1", x"ff1", x"ff1", x"ff0", x"ff0",
        x"ff0", x"fef", x"fef", x"fee", x"fee", x"fee", x"fed", x"fed",
        x"fec", x"fec", x"fec", x"feb", x"feb", x"fea", x"fea", x"fe9",
        x"fe9", x"fe8", x"fe8", x"fe7", x"fe7", x"fe6", x"fe6", x"fe5",
        x"fe5", x"fe4", x"fe4", x"fe3", x"fe3", x"fe2", x"fe2", x"fe1",
        x"fe1", x"fe0", x"fe0", x"fdf", x"fdf", x"fde", x"fde", x"fdd",
        x"fdc", x"fdc", x"fdb", x"fdb", x"fda", x"fd9", x"fd9", x"fd8",
        x"fd8", x"fd7", x"fd6", x"fd6", x"fd5", x"fd5", x"fd4", x"fd3",
        x"fd3", x"fd2", x"fd1", x"fd1", x"fd0", x"fcf", x"fcf", x"fce",
        x"fcd", x"fcd", x"fcc", x"fcb", x"fca", x"fca", x"fc9", x"fc8",
        x"fc8", x"fc7", x"fc6", x"fc5", x"fc5", x"fc4", x"fc3", x"fc2",
        x"fc2", x"fc1", x"fc0", x"fbf", x"fbf", x"fbe", x"fbd", x"fbc",
        x"fbb", x"fbb", x"fba", x"fb9", x"fb8", x"fb7", x"fb6", x"fb6",
        x"fb5", x"fb4", x"fb3", x"fb2", x"fb1", x"fb1", x"fb0", x"faf",
        x"fae", x"fad", x"fac", x"fab", x"faa", x"faa", x"fa9", x"fa8",
        x"fa7", x"fa6", x"fa5", x"fa4", x"fa3", x"fa2", x"fa1", x"fa0",
        x"f9f", x"f9e", x"f9d", x"f9d", x"f9c", x"f9b", x"f9a", x"f99",
        x"f98", x"f97", x"f96", x"f95", x"f94", x"f93", x"f92", x"f91",
        x"f90", x"f8f", x"f8e", x"f8d", x"f8c", x"f8a", x"f89", x"f88",
        x"f87", x"f86", x"f85", x"f84", x"f83", x"f82", x"f81", x"f80",
        x"f7f", x"f7e", x"f7d", x"f7b", x"f7a", x"f79", x"f78", x"f77",
        x"f76", x"f75", x"f74", x"f72", x"f71", x"f70", x"f6f", x"f6e",
        x"f6d", x"f6b", x"f6a", x"f69", x"f68", x"f67", x"f66", x"f64",
        x"f63", x"f62", x"f61", x"f60", x"f5e", x"f5d", x"f5c", x"f5b",
        x"f59", x"f58", x"f57", x"f56", x"f54", x"f53", x"f52", x"f51",
        x"f4f", x"f4e", x"f4d", x"f4c", x"f4a", x"f49", x"f48", x"f46",
        x"f45", x"f44", x"f42", x"f41", x"f40", x"f3e", x"f3d", x"f3c",
        x"f3a", x"f39", x"f38", x"f36", x"f35", x"f34", x"f32", x"f31",
        x"f30", x"f2e", x"f2d", x"f2b", x"f2a", x"f29", x"f27", x"f26",
        x"f24", x"f23", x"f22", x"f20", x"f1f", x"f1d", x"f1c", x"f1a",
        x"f19", x"f17", x"f16", x"f15", x"f13", x"f12", x"f10", x"f0f",
        x"f0d", x"f0c", x"f0a", x"f09", x"f07", x"f06", x"f04", x"f03",
        x"f01", x"f00", x"efe", x"efd", x"efb", x"efa", x"ef8", x"ef7",
        x"ef5", x"ef3", x"ef2", x"ef0", x"eef", x"eed", x"eec", x"eea",
        x"ee8", x"ee7", x"ee5", x"ee4", x"ee2", x"ee1", x"edf", x"edd",
        x"edc", x"eda", x"ed8", x"ed7", x"ed5", x"ed4", x"ed2", x"ed0",
        x"ecf", x"ecd", x"ecb", x"eca", x"ec8", x"ec6", x"ec5", x"ec3",
        x"ec1", x"ec0", x"ebe", x"ebc", x"ebb", x"eb9", x"eb7", x"eb5",
        x"eb4", x"eb2", x"eb0", x"eaf", x"ead", x"eab", x"ea9", x"ea8",
        x"ea6", x"ea4", x"ea2", x"ea1", x"e9f", x"e9d", x"e9b", x"e9a",
        x"e98", x"e96", x"e94", x"e92", x"e91", x"e8f", x"e8d", x"e8b",
        x"e8a", x"e88", x"e86", x"e84", x"e82", x"e80", x"e7f", x"e7d",
        x"e7b", x"e79", x"e77", x"e75", x"e74", x"e72", x"e70", x"e6e",
        x"e6c", x"e6a", x"e68", x"e66", x"e65", x"e63", x"e61", x"e5f",
        x"e5d", x"e5b", x"e59", x"e57", x"e55", x"e53", x"e51", x"e50",
        x"e4e", x"e4c", x"e4a", x"e48", x"e46", x"e44", x"e42", x"e40",
        x"e3e", x"e3c", x"e3a", x"e38", x"e36", x"e34", x"e32", x"e30",
        x"e2e", x"e2c", x"e2a", x"e28", x"e26", x"e24", x"e22", x"e20",
        x"e1e", x"e1c", x"e1a", x"e18", x"e16", x"e14", x"e12", x"e10",
        x"e0e", x"e0c", x"e0a", x"e08", x"e06", x"e04", x"e02", x"dff",
        x"dfd", x"dfb", x"df9", x"df7", x"df5", x"df3", x"df1", x"def",
        x"ded", x"dea", x"de8", x"de6", x"de4", x"de2", x"de0", x"dde",
        x"ddc", x"dd9", x"dd7", x"dd5", x"dd3", x"dd1", x"dcf", x"dcd",
        x"dca", x"dc8", x"dc6", x"dc4", x"dc2", x"dc0", x"dbd", x"dbb",
        x"db9", x"db7", x"db5", x"db2", x"db0", x"dae", x"dac", x"daa",
        x"da7", x"da5", x"da3", x"da1", x"d9e", x"d9c", x"d9a", x"d98",
        x"d95", x"d93", x"d91", x"d8f", x"d8c", x"d8a", x"d88", x"d86",
        x"d83", x"d81", x"d7f", x"d7c", x"d7a", x"d78", x"d76", x"d73",
        x"d71", x"d6f", x"d6c", x"d6a", x"d68", x"d65", x"d63", x"d61",
        x"d5f", x"d5c", x"d5a", x"d58", x"d55", x"d53", x"d50", x"d4e",
        x"d4c", x"d49", x"d47", x"d45", x"d42", x"d40", x"d3e", x"d3b",
        x"d39", x"d36", x"d34", x"d32", x"d2f", x"d2d", x"d2b", x"d28",
        x"d26", x"d23", x"d21", x"d1f", x"d1c", x"d1a", x"d17", x"d15",
        x"d12", x"d10", x"d0e", x"d0b", x"d09", x"d06", x"d04", x"d01",
        x"cff", x"cfc", x"cfa", x"cf8", x"cf5", x"cf3", x"cf0", x"cee",
        x"ceb", x"ce9", x"ce6", x"ce4", x"ce1", x"cdf", x"cdc", x"cda",
        x"cd7", x"cd5", x"cd2", x"cd0", x"ccd", x"ccb", x"cc8", x"cc6",
        x"cc3", x"cc1", x"cbe", x"cbc", x"cb9", x"cb7", x"cb4", x"cb1",
        x"caf", x"cac", x"caa", x"ca7", x"ca5", x"ca2", x"ca0", x"c9d",
        x"c9a", x"c98", x"c95", x"c93", x"c90", x"c8e", x"c8b", x"c88",
        x"c86", x"c83", x"c81", x"c7e", x"c7b", x"c79", x"c76", x"c74",
        x"c71", x"c6e", x"c6c", x"c69", x"c67", x"c64", x"c61", x"c5f",
        x"c5c", x"c59", x"c57", x"c54", x"c52", x"c4f", x"c4c", x"c4a",
        x"c47", x"c44", x"c42", x"c3f", x"c3c", x"c3a", x"c37", x"c34",
        x"c32", x"c2f", x"c2c", x"c2a", x"c27", x"c24", x"c22", x"c1f",
        x"c1c", x"c19", x"c17", x"c14", x"c11", x"c0f", x"c0c", x"c09",
        x"c06", x"c04", x"c01", x"bfe", x"bfc", x"bf9", x"bf6", x"bf3",
        x"bf1", x"bee", x"beb", x"be9", x"be6", x"be3", x"be0", x"bde",
        x"bdb", x"bd8", x"bd5", x"bd3", x"bd0", x"bcd", x"bca", x"bc7",
        x"bc5", x"bc2", x"bbf", x"bbc", x"bba", x"bb7", x"bb4", x"bb1",
        x"bae", x"bac", x"ba9", x"ba6", x"ba3", x"ba0", x"b9e", x"b9b",
        x"b98", x"b95", x"b92", x"b90", x"b8d", x"b8a", x"b87", x"b84",
        x"b82", x"b7f", x"b7c", x"b79", x"b76", x"b73", x"b71", x"b6e",
        x"b6b", x"b68", x"b65", x"b62", x"b60", x"b5d", x"b5a", x"b57",
        x"b54", x"b51", x"b4e", x"b4c", x"b49", x"b46", x"b43", x"b40",
        x"b3d", x"b3a", x"b37", x"b35", x"b32", x"b2f", x"b2c", x"b29",
        x"b26", x"b23", x"b20", x"b1e", x"b1b", x"b18", x"b15", x"b12",
        x"b0f", x"b0c", x"b09", x"b06", x"b03", x"b01", x"afe", x"afb",
        x"af8", x"af5", x"af2", x"aef", x"aec", x"ae9", x"ae6", x"ae3",
        x"ae0", x"add", x"adb", x"ad8", x"ad5", x"ad2", x"acf", x"acc",
        x"ac9", x"ac6", x"ac3", x"ac0", x"abd", x"aba", x"ab7", x"ab4",
        x"ab1", x"aae", x"aab", x"aa8", x"aa5", x"aa2", x"aa0", x"a9d",
        x"a9a", x"a97", x"a94", x"a91", x"a8e", x"a8b", x"a88", x"a85",
        x"a82", x"a7f", x"a7c", x"a79", x"a76", x"a73", x"a70", x"a6d",
        x"a6a", x"a67", x"a64", x"a61", x"a5e", x"a5b", x"a58", x"a55",
        x"a52", x"a4f", x"a4c", x"a49", x"a46", x"a43", x"a40", x"a3d",
        x"a3a", x"a37", x"a34", x"a31", x"a2e", x"a2b", x"a28", x"a25",
        x"a22", x"a1f", x"a1c", x"a19", x"a15", x"a12", x"a0f", x"a0c",
        x"a09", x"a06", x"a03", x"a00", x"9fd", x"9fa", x"9f7", x"9f4",
        x"9f1", x"9ee", x"9eb", x"9e8", x"9e5", x"9e2", x"9df", x"9dc",
        x"9d9", x"9d6", x"9d2", x"9cf", x"9cc", x"9c9", x"9c6", x"9c3",
        x"9c0", x"9bd", x"9ba", x"9b7", x"9b4", x"9b1", x"9ae", x"9ab",
        x"9a8", x"9a4", x"9a1", x"99e", x"99b", x"998", x"995", x"992",
        x"98f", x"98c", x"989", x"986", x"983", x"980", x"97c", x"979",
        x"976", x"973", x"970", x"96d", x"96a", x"967", x"964", x"961",
        x"95e", x"95a", x"957", x"954", x"951", x"94e", x"94b", x"948",
        x"945", x"942", x"93f", x"93b", x"938", x"935", x"932", x"92f",
        x"92c", x"929", x"926", x"923", x"91f", x"91c", x"919", x"916",
        x"913", x"910", x"90d", x"90a", x"907", x"903", x"900", x"8fd",
        x"8fa", x"8f7", x"8f4", x"8f1", x"8ee", x"8eb", x"8e7", x"8e4",
        x"8e1", x"8de", x"8db", x"8d8", x"8d5", x"8d2", x"8ce", x"8cb",
        x"8c8", x"8c5", x"8c2", x"8bf", x"8bc", x"8b9", x"8b5", x"8b2",
        x"8af", x"8ac", x"8a9", x"8a6", x"8a3", x"8a0", x"89c", x"899",
        x"896", x"893", x"890", x"88d", x"88a", x"886", x"883", x"880",
        x"87d", x"87a", x"877", x"874", x"871", x"86d", x"86a", x"867",
        x"864", x"861", x"85e", x"85b", x"857", x"854", x"851", x"84e",
        x"84b", x"848", x"845", x"841", x"83e", x"83b", x"838", x"835",
        x"832", x"82f", x"82b", x"828", x"825", x"822", x"81f", x"81c",
        x"819", x"815", x"812", x"80f", x"80c", x"809", x"806", x"803",
        x"800", x"7fc", x"7f9", x"7f6", x"7f3", x"7f0", x"7ed", x"7ea",
        x"7e6", x"7e3", x"7e0", x"7dd", x"7da", x"7d7", x"7d4", x"7d0",
        x"7cd", x"7ca", x"7c7", x"7c4", x"7c1", x"7be", x"7ba", x"7b7",
        x"7b4", x"7b1", x"7ae", x"7ab", x"7a8", x"7a4", x"7a1", x"79e",
        x"79b", x"798", x"795", x"792", x"78e", x"78b", x"788", x"785",
        x"782", x"77f", x"77c", x"779", x"775", x"772", x"76f", x"76c",
        x"769", x"766", x"763", x"75f", x"75c", x"759", x"756", x"753",
        x"750", x"74d", x"74a", x"746", x"743", x"740", x"73d", x"73a",
        x"737", x"734", x"731", x"72d", x"72a", x"727", x"724", x"721",
        x"71e", x"71b", x"718", x"714", x"711", x"70e", x"70b", x"708",
        x"705", x"702", x"6ff", x"6fc", x"6f8", x"6f5", x"6f2", x"6ef",
        x"6ec", x"6e9", x"6e6", x"6e3", x"6e0", x"6dc", x"6d9", x"6d6",
        x"6d3", x"6d0", x"6cd", x"6ca", x"6c7", x"6c4", x"6c0", x"6bd",
        x"6ba", x"6b7", x"6b4", x"6b1", x"6ae", x"6ab", x"6a8", x"6a5",
        x"6a1", x"69e", x"69b", x"698", x"695", x"692", x"68f", x"68c",
        x"689", x"686", x"683", x"67f", x"67c", x"679", x"676", x"673",
        x"670", x"66d", x"66a", x"667", x"664", x"661", x"65e", x"65b",
        x"657", x"654", x"651", x"64e", x"64b", x"648", x"645", x"642",
        x"63f", x"63c", x"639", x"636", x"633", x"630", x"62d", x"629",
        x"626", x"623", x"620", x"61d", x"61a", x"617", x"614", x"611",
        x"60e", x"60b", x"608", x"605", x"602", x"5ff", x"5fc", x"5f9",
        x"5f6", x"5f3", x"5f0", x"5ed", x"5ea", x"5e6", x"5e3", x"5e0",
        x"5dd", x"5da", x"5d7", x"5d4", x"5d1", x"5ce", x"5cb", x"5c8",
        x"5c5", x"5c2", x"5bf", x"5bc", x"5b9", x"5b6", x"5b3", x"5b0",
        x"5ad", x"5aa", x"5a7", x"5a4", x"5a1", x"59e", x"59b", x"598",
        x"595", x"592", x"58f", x"58c", x"589", x"586", x"583", x"580",
        x"57d", x"57a", x"577", x"574", x"571", x"56e", x"56b", x"568",
        x"565", x"562", x"55f", x"55d", x"55a", x"557", x"554", x"551",
        x"54e", x"54b", x"548", x"545", x"542", x"53f", x"53c", x"539",
        x"536", x"533", x"530", x"52d", x"52a", x"527", x"524", x"522",
        x"51f", x"51c", x"519", x"516", x"513", x"510", x"50d", x"50a",
        x"507", x"504", x"501", x"4fe", x"4fc", x"4f9", x"4f6", x"4f3",
        x"4f0", x"4ed", x"4ea", x"4e7", x"4e4", x"4e1", x"4df", x"4dc",
        x"4d9", x"4d6", x"4d3", x"4d0", x"4cd", x"4ca", x"4c8", x"4c5",
        x"4c2", x"4bf", x"4bc", x"4b9", x"4b6", x"4b3", x"4b1", x"4ae",
        x"4ab", x"4a8", x"4a5", x"4a2", x"49f", x"49d", x"49a", x"497",
        x"494", x"491", x"48e", x"48c", x"489", x"486", x"483", x"480",
        x"47d", x"47b", x"478", x"475", x"472", x"46f", x"46d", x"46a",
        x"467", x"464", x"461", x"45f", x"45c", x"459", x"456", x"453",
        x"451", x"44e", x"44b", x"448", x"445", x"443", x"440", x"43d",
        x"43a", x"438", x"435", x"432", x"42f", x"42c", x"42a", x"427",
        x"424", x"421", x"41f", x"41c", x"419", x"416", x"414", x"411",
        x"40e", x"40c", x"409", x"406", x"403", x"401", x"3fe", x"3fb",
        x"3f9", x"3f6", x"3f3", x"3f0", x"3ee", x"3eb", x"3e8", x"3e6",
        x"3e3", x"3e0", x"3dd", x"3db", x"3d8", x"3d5", x"3d3", x"3d0",
        x"3cd", x"3cb", x"3c8", x"3c5", x"3c3", x"3c0", x"3bd", x"3bb",
        x"3b8", x"3b5", x"3b3", x"3b0", x"3ad", x"3ab", x"3a8", x"3a6",
        x"3a3", x"3a0", x"39e", x"39b", x"398", x"396", x"393", x"391",
        x"38e", x"38b", x"389", x"386", x"384", x"381", x"37e", x"37c",
        x"379", x"377", x"374", x"371", x"36f", x"36c", x"36a", x"367",
        x"365", x"362", x"35f", x"35d", x"35a", x"358", x"355", x"353",
        x"350", x"34e", x"34b", x"348", x"346", x"343", x"341", x"33e",
        x"33c", x"339", x"337", x"334", x"332", x"32f", x"32d", x"32a",
        x"328", x"325", x"323", x"320", x"31e", x"31b", x"319", x"316",
        x"314", x"311", x"30f", x"30c", x"30a", x"307", x"305", x"303",
        x"300", x"2fe", x"2fb", x"2f9", x"2f6", x"2f4", x"2f1", x"2ef",
        x"2ed", x"2ea", x"2e8", x"2e5", x"2e3", x"2e0", x"2de", x"2dc",
        x"2d9", x"2d7", x"2d4", x"2d2", x"2d0", x"2cd", x"2cb", x"2c9",
        x"2c6", x"2c4", x"2c1", x"2bf", x"2bd", x"2ba", x"2b8", x"2b6",
        x"2b3", x"2b1", x"2af", x"2ac", x"2aa", x"2a7", x"2a5", x"2a3",
        x"2a0", x"29e", x"29c", x"29a", x"297", x"295", x"293", x"290",
        x"28e", x"28c", x"289", x"287", x"285", x"283", x"280", x"27e",
        x"27c", x"279", x"277", x"275", x"273", x"270", x"26e", x"26c",
        x"26a", x"267", x"265", x"263", x"261", x"25e", x"25c", x"25a",
        x"258", x"255", x"253", x"251", x"24f", x"24d", x"24a", x"248",
        x"246", x"244", x"242", x"23f", x"23d", x"23b", x"239", x"237",
        x"235", x"232", x"230", x"22e", x"22c", x"22a", x"228", x"226",
        x"223", x"221", x"21f", x"21d", x"21b", x"219", x"217", x"215",
        x"212", x"210", x"20e", x"20c", x"20a", x"208", x"206", x"204",
        x"202", x"200", x"1fd", x"1fb", x"1f9", x"1f7", x"1f5", x"1f3",
        x"1f1", x"1ef", x"1ed", x"1eb", x"1e9", x"1e7", x"1e5", x"1e3",
        x"1e1", x"1df", x"1dd", x"1db", x"1d9", x"1d7", x"1d5", x"1d3",
        x"1d1", x"1cf", x"1cd", x"1cb", x"1c9", x"1c7", x"1c5", x"1c3",
        x"1c1", x"1bf", x"1bd", x"1bb", x"1b9", x"1b7", x"1b5", x"1b3",
        x"1b1", x"1af", x"1ae", x"1ac", x"1aa", x"1a8", x"1a6", x"1a4",
        x"1a2", x"1a0", x"19e", x"19c", x"19a", x"199", x"197", x"195",
        x"193", x"191", x"18f", x"18d", x"18b", x"18a", x"188", x"186",
        x"184", x"182", x"180", x"17f", x"17d", x"17b", x"179", x"177",
        x"175", x"174", x"172", x"170", x"16e", x"16d", x"16b", x"169",
        x"167", x"165", x"164", x"162", x"160", x"15e", x"15d", x"15b",
        x"159", x"157", x"156", x"154", x"152", x"150", x"14f", x"14d",
        x"14b", x"14a", x"148", x"146", x"144", x"143", x"141", x"13f",
        x"13e", x"13c", x"13a", x"139", x"137", x"135", x"134", x"132",
        x"130", x"12f", x"12d", x"12b", x"12a", x"128", x"127", x"125",
        x"123", x"122", x"120", x"11e", x"11d", x"11b", x"11a", x"118",
        x"117", x"115", x"113", x"112", x"110", x"10f", x"10d", x"10c",
        x"10a", x"108", x"107", x"105", x"104", x"102", x"101", x"0ff",
        x"0fe", x"0fc", x"0fb", x"0f9", x"0f8", x"0f6", x"0f5", x"0f3",
        x"0f2", x"0f0", x"0ef", x"0ed", x"0ec", x"0ea", x"0e9", x"0e8",
        x"0e6", x"0e5", x"0e3", x"0e2", x"0e0", x"0df", x"0dd", x"0dc",
        x"0db", x"0d9", x"0d8", x"0d6", x"0d5", x"0d4", x"0d2", x"0d1",
        x"0cf", x"0ce", x"0cd", x"0cb", x"0ca", x"0c9", x"0c7", x"0c6",
        x"0c5", x"0c3", x"0c2", x"0c1", x"0bf", x"0be", x"0bd", x"0bb",
        x"0ba", x"0b9", x"0b7", x"0b6", x"0b5", x"0b3", x"0b2", x"0b1",
        x"0b0", x"0ae", x"0ad", x"0ac", x"0ab", x"0a9", x"0a8", x"0a7",
        x"0a6", x"0a4", x"0a3", x"0a2", x"0a1", x"09f", x"09e", x"09d",
        x"09c", x"09b", x"099", x"098", x"097", x"096", x"095", x"094",
        x"092", x"091", x"090", x"08f", x"08e", x"08d", x"08b", x"08a",
        x"089", x"088", x"087", x"086", x"085", x"084", x"082", x"081",
        x"080", x"07f", x"07e", x"07d", x"07c", x"07b", x"07a", x"079",
        x"078", x"077", x"076", x"075", x"073", x"072", x"071", x"070",
        x"06f", x"06e", x"06d", x"06c", x"06b", x"06a", x"069", x"068",
        x"067", x"066", x"065", x"064", x"063", x"062", x"062", x"061",
        x"060", x"05f", x"05e", x"05d", x"05c", x"05b", x"05a", x"059",
        x"058", x"057", x"056", x"055", x"055", x"054", x"053", x"052",
        x"051", x"050", x"04f", x"04e", x"04e", x"04d", x"04c", x"04b",
        x"04a", x"049", x"049", x"048", x"047", x"046", x"045", x"044",
        x"044", x"043", x"042", x"041", x"040", x"040", x"03f", x"03e",
        x"03d", x"03d", x"03c", x"03b", x"03a", x"03a", x"039", x"038",
        x"037", x"037", x"036", x"035", x"035", x"034", x"033", x"032",
        x"032", x"031", x"030", x"030", x"02f", x"02e", x"02e", x"02d",
        x"02c", x"02c", x"02b", x"02a", x"02a", x"029", x"029", x"028",
        x"027", x"027", x"026", x"026", x"025", x"024", x"024", x"023",
        x"023", x"022", x"021", x"021", x"020", x"020", x"01f", x"01f",
        x"01e", x"01e", x"01d", x"01d", x"01c", x"01c", x"01b", x"01b",
        x"01a", x"01a", x"019", x"019", x"018", x"018", x"017", x"017",
        x"016", x"016", x"015", x"015", x"014", x"014", x"013", x"013",
        x"013", x"012", x"012", x"011", x"011", x"011", x"010", x"010",
        x"00f", x"00f", x"00f", x"00e", x"00e", x"00e", x"00d", x"00d",
        x"00c", x"00c", x"00c", x"00b", x"00b", x"00b", x"00a", x"00a",
        x"00a", x"00a", x"009", x"009", x"009", x"008", x"008", x"008",
        x"008", x"007", x"007", x"007", x"007", x"006", x"006", x"006",
        x"006", x"005", x"005", x"005", x"005", x"004", x"004", x"004",
        x"004", x"004", x"003", x"003", x"003", x"003", x"003", x"003",
        x"002", x"002", x"002", x"002", x"002", x"002", x"002", x"002",
        x"001", x"001", x"001", x"001", x"001", x"001", x"001", x"001",
        x"001", x"001", x"000", x"000", x"000", x"000", x"000", x"000",
        x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
        x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
        x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"001",
        x"001", x"001", x"001", x"001", x"001", x"001", x"001", x"001",
        x"001", x"002", x"002", x"002", x"002", x"002", x"002", x"002",
        x"002", x"003", x"003", x"003", x"003", x"003", x"003", x"004",
        x"004", x"004", x"004", x"004", x"005", x"005", x"005", x"005",
        x"006", x"006", x"006", x"006", x"007", x"007", x"007", x"007",
        x"008", x"008", x"008", x"008", x"009", x"009", x"009", x"00a",
        x"00a", x"00a", x"00a", x"00b", x"00b", x"00b", x"00c", x"00c",
        x"00c", x"00d", x"00d", x"00e", x"00e", x"00e", x"00f", x"00f",
        x"00f", x"010", x"010", x"011", x"011", x"011", x"012", x"012",
        x"013", x"013", x"013", x"014", x"014", x"015", x"015", x"016",
        x"016", x"017", x"017", x"018", x"018", x"019", x"019", x"01a",
        x"01a", x"01b", x"01b", x"01c", x"01c", x"01d", x"01d", x"01e",
        x"01e", x"01f", x"01f", x"020", x"020", x"021", x"021", x"022",
        x"023", x"023", x"024", x"024", x"025", x"026", x"026", x"027",
        x"027", x"028", x"029", x"029", x"02a", x"02a", x"02b", x"02c",
        x"02c", x"02d", x"02e", x"02e", x"02f", x"030", x"030", x"031",
        x"032", x"032", x"033", x"034", x"035", x"035", x"036", x"037",
        x"037", x"038", x"039", x"03a", x"03a", x"03b", x"03c", x"03d",
        x"03d", x"03e", x"03f", x"040", x"040", x"041", x"042", x"043",
        x"044", x"044", x"045", x"046", x"047", x"048", x"049", x"049",
        x"04a", x"04b", x"04c", x"04d", x"04e", x"04e", x"04f", x"050",
        x"051", x"052", x"053", x"054", x"055", x"055", x"056", x"057",
        x"058", x"059", x"05a", x"05b", x"05c", x"05d", x"05e", x"05f",
        x"060", x"061", x"062", x"062", x"063", x"064", x"065", x"066",
        x"067", x"068", x"069", x"06a", x"06b", x"06c", x"06d", x"06e",
        x"06f", x"070", x"071", x"072", x"073", x"075", x"076", x"077",
        x"078", x"079", x"07a", x"07b", x"07c", x"07d", x"07e", x"07f",
        x"080", x"081", x"082", x"084", x"085", x"086", x"087", x"088",
        x"089", x"08a", x"08b", x"08d", x"08e", x"08f", x"090", x"091",
        x"092", x"094", x"095", x"096", x"097", x"098", x"099", x"09b",
        x"09c", x"09d", x"09e", x"09f", x"0a1", x"0a2", x"0a3", x"0a4",
        x"0a6", x"0a7", x"0a8", x"0a9", x"0ab", x"0ac", x"0ad", x"0ae",
        x"0b0", x"0b1", x"0b2", x"0b3", x"0b5", x"0b6", x"0b7", x"0b9",
        x"0ba", x"0bb", x"0bd", x"0be", x"0bf", x"0c1", x"0c2", x"0c3",
        x"0c5", x"0c6", x"0c7", x"0c9", x"0ca", x"0cb", x"0cd", x"0ce",
        x"0cf", x"0d1", x"0d2", x"0d4", x"0d5", x"0d6", x"0d8", x"0d9",
        x"0db", x"0dc", x"0dd", x"0df", x"0e0", x"0e2", x"0e3", x"0e5",
        x"0e6", x"0e8", x"0e9", x"0ea", x"0ec", x"0ed", x"0ef", x"0f0",
        x"0f2", x"0f3", x"0f5", x"0f6", x"0f8", x"0f9", x"0fb", x"0fc",
        x"0fe", x"0ff", x"101", x"102", x"104", x"105", x"107", x"108",
        x"10a", x"10c", x"10d", x"10f", x"110", x"112", x"113", x"115",
        x"117", x"118", x"11a", x"11b", x"11d", x"11e", x"120", x"122",
        x"123", x"125", x"127", x"128", x"12a", x"12b", x"12d", x"12f",
        x"130", x"132", x"134", x"135", x"137", x"139", x"13a", x"13c",
        x"13e", x"13f", x"141", x"143", x"144", x"146", x"148", x"14a",
        x"14b", x"14d", x"14f", x"150", x"152", x"154", x"156", x"157",
        x"159", x"15b", x"15d", x"15e", x"160", x"162", x"164", x"165",
        x"167", x"169", x"16b", x"16d", x"16e", x"170", x"172", x"174",
        x"175", x"177", x"179", x"17b", x"17d", x"17f", x"180", x"182",
        x"184", x"186", x"188", x"18a", x"18b", x"18d", x"18f", x"191",
        x"193", x"195", x"197", x"199", x"19a", x"19c", x"19e", x"1a0",
        x"1a2", x"1a4", x"1a6", x"1a8", x"1aa", x"1ac", x"1ae", x"1af",
        x"1b1", x"1b3", x"1b5", x"1b7", x"1b9", x"1bb", x"1bd", x"1bf",
        x"1c1", x"1c3", x"1c5", x"1c7", x"1c9", x"1cb", x"1cd", x"1cf",
        x"1d1", x"1d3", x"1d5", x"1d7", x"1d9", x"1db", x"1dd", x"1df",
        x"1e1", x"1e3", x"1e5", x"1e7", x"1e9", x"1eb", x"1ed", x"1ef",
        x"1f1", x"1f3", x"1f5", x"1f7", x"1f9", x"1fb", x"1fd", x"200",
        x"202", x"204", x"206", x"208", x"20a", x"20c", x"20e", x"210",
        x"212", x"215", x"217", x"219", x"21b", x"21d", x"21f", x"221",
        x"223", x"226", x"228", x"22a", x"22c", x"22e", x"230", x"232",
        x"235", x"237", x"239", x"23b", x"23d", x"23f", x"242", x"244",
        x"246", x"248", x"24a", x"24d", x"24f", x"251", x"253", x"255",
        x"258", x"25a", x"25c", x"25e", x"261", x"263", x"265", x"267",
        x"26a", x"26c", x"26e", x"270", x"273", x"275", x"277", x"279",
        x"27c", x"27e", x"280", x"283", x"285", x"287", x"289", x"28c",
        x"28e", x"290", x"293", x"295", x"297", x"29a", x"29c", x"29e",
        x"2a0", x"2a3", x"2a5", x"2a7", x"2aa", x"2ac", x"2af", x"2b1",
        x"2b3", x"2b6", x"2b8", x"2ba", x"2bd", x"2bf", x"2c1", x"2c4",
        x"2c6", x"2c9", x"2cb", x"2cd", x"2d0", x"2d2", x"2d4", x"2d7",
        x"2d9", x"2dc", x"2de", x"2e0", x"2e3", x"2e5", x"2e8", x"2ea",
        x"2ed", x"2ef", x"2f1", x"2f4", x"2f6", x"2f9", x"2fb", x"2fe",
        x"300", x"303", x"305", x"307", x"30a", x"30c", x"30f", x"311",
        x"314", x"316", x"319", x"31b", x"31e", x"320", x"323", x"325",
        x"328", x"32a", x"32d", x"32f", x"332", x"334", x"337", x"339",
        x"33c", x"33e", x"341", x"343", x"346", x"348", x"34b", x"34e",
        x"350", x"353", x"355", x"358", x"35a", x"35d", x"35f", x"362",
        x"365", x"367", x"36a", x"36c", x"36f", x"371", x"374", x"377",
        x"379", x"37c", x"37e", x"381", x"384", x"386", x"389", x"38b",
        x"38e", x"391", x"393", x"396", x"398", x"39b", x"39e", x"3a0",
        x"3a3", x"3a6", x"3a8", x"3ab", x"3ad", x"3b0", x"3b3", x"3b5",
        x"3b8", x"3bb", x"3bd", x"3c0", x"3c3", x"3c5", x"3c8", x"3cb",
        x"3cd", x"3d0", x"3d3", x"3d5", x"3d8", x"3db", x"3dd", x"3e0",
        x"3e3", x"3e6", x"3e8", x"3eb", x"3ee", x"3f0", x"3f3", x"3f6",
        x"3f9", x"3fb", x"3fe", x"401", x"403", x"406", x"409", x"40c",
        x"40e", x"411", x"414", x"416", x"419", x"41c", x"41f", x"421",
        x"424", x"427", x"42a", x"42c", x"42f", x"432", x"435", x"438",
        x"43a", x"43d", x"440", x"443", x"445", x"448", x"44b", x"44e",
        x"451", x"453", x"456", x"459", x"45c", x"45f", x"461", x"464",
        x"467", x"46a", x"46d", x"46f", x"472", x"475", x"478", x"47b",
        x"47d", x"480", x"483", x"486", x"489", x"48c", x"48e", x"491",
        x"494", x"497", x"49a", x"49d", x"49f", x"4a2", x"4a5", x"4a8",
        x"4ab", x"4ae", x"4b1", x"4b3", x"4b6", x"4b9", x"4bc", x"4bf",
        x"4c2", x"4c5", x"4c8", x"4ca", x"4cd", x"4d0", x"4d3", x"4d6",
        x"4d9", x"4dc", x"4df", x"4e1", x"4e4", x"4e7", x"4ea", x"4ed",
        x"4f0", x"4f3", x"4f6", x"4f9", x"4fc", x"4fe", x"501", x"504",
        x"507", x"50a", x"50d", x"510", x"513", x"516", x"519", x"51c",
        x"51f", x"522", x"524", x"527", x"52a", x"52d", x"530", x"533",
        x"536", x"539", x"53c", x"53f", x"542", x"545", x"548", x"54b",
        x"54e", x"551", x"554", x"557", x"55a", x"55d", x"55f", x"562",
        x"565", x"568", x"56b", x"56e", x"571", x"574", x"577", x"57a",
        x"57d", x"580", x"583", x"586", x"589", x"58c", x"58f", x"592",
        x"595", x"598", x"59b", x"59e", x"5a1", x"5a4", x"5a7", x"5aa",
        x"5ad", x"5b0", x"5b3", x"5b6", x"5b9", x"5bc", x"5bf", x"5c2",
        x"5c5", x"5c8", x"5cb", x"5ce", x"5d1", x"5d4", x"5d7", x"5da",
        x"5dd", x"5e0", x"5e3", x"5e6", x"5ea", x"5ed", x"5f0", x"5f3",
        x"5f6", x"5f9", x"5fc", x"5ff", x"602", x"605", x"608", x"60b",
        x"60e", x"611", x"614", x"617", x"61a", x"61d", x"620", x"623",
        x"626", x"629", x"62d", x"630", x"633", x"636", x"639", x"63c",
        x"63f", x"642", x"645", x"648", x"64b", x"64e", x"651", x"654",
        x"657", x"65b", x"65e", x"661", x"664", x"667", x"66a", x"66d",
        x"670", x"673", x"676", x"679", x"67c", x"67f", x"683", x"686",
        x"689", x"68c", x"68f", x"692", x"695", x"698", x"69b", x"69e",
        x"6a1", x"6a5", x"6a8", x"6ab", x"6ae", x"6b1", x"6b4", x"6b7",
        x"6ba", x"6bd", x"6c0", x"6c4", x"6c7", x"6ca", x"6cd", x"6d0",
        x"6d3", x"6d6", x"6d9", x"6dc", x"6e0", x"6e3", x"6e6", x"6e9",
        x"6ec", x"6ef", x"6f2", x"6f5", x"6f8", x"6fc", x"6ff", x"702",
        x"705", x"708", x"70b", x"70e", x"711", x"714", x"718", x"71b",
        x"71e", x"721", x"724", x"727", x"72a", x"72d", x"731", x"734",
        x"737", x"73a", x"73d", x"740", x"743", x"746", x"74a", x"74d",
        x"750", x"753", x"756", x"759", x"75c", x"75f", x"763", x"766",
        x"769", x"76c", x"76f", x"772", x"775", x"779", x"77c", x"77f",
        x"782", x"785", x"788", x"78b", x"78e", x"792", x"795", x"798",
        x"79b", x"79e", x"7a1", x"7a4", x"7a8", x"7ab", x"7ae", x"7b1",
        x"7b4", x"7b7", x"7ba", x"7be", x"7c1", x"7c4", x"7c7", x"7ca",
        x"7cd", x"7d0", x"7d4", x"7d7", x"7da", x"7dd", x"7e0", x"7e3",
        x"7e6", x"7ea", x"7ed", x"7f0", x"7f3", x"7f6", x"7f9", x"7fc"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr,clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp,en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
