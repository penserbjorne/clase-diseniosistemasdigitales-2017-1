library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity rom_vicflo is
    port (
        clk  : in  std_logic;
        en   : in  std_logic := '1';
        addr : in  std_logic_vector(10 downto 0);
        data : out std_logic_vector(11 downto 0)
    );
end rom_vicflo;

architecture arch of rom_vicflo is
    type memoria_rom is array (0 to 2047) of std_logic_vector (11 downto 0);
    constant ROM : memoria_rom := (
        x"7f9", x"7ed", x"7e0", x"7d3", x"7c7", x"7ba", x"7ae", x"7a1",
        x"795", x"788", x"77c", x"76f", x"762", x"756", x"749", x"73d", 
        x"730", x"724", x"717", x"70b", x"6fe", x"6f2", x"6e5", x"6d9",
        x"6cd", x"6c0", x"6b4", x"6a7", x"69b", x"68f", x"682", x"676",
        x"66a", x"65d", x"651", x"645", x"638", x"62c", x"620", x"614",
        x"607", x"5fb", x"5ef", x"5e3", x"5d7", x"5cb", x"5bf", x"5b3",
        x"5a7", x"59b", x"58f", x"583", x"577", x"56b", x"55f", x"553",
        x"547", x"53b", x"530", x"524", x"518", x"50c", x"501", x"4f5",
        x"4e9", x"4de", x"4d2", x"4c7", x"4bb", x"4b0", x"4a4", x"499",
        x"48e", x"482", x"477", x"46c", x"460", x"455", x"44a", x"43f",
        x"434", x"429", x"41e", x"413", x"408", x"3fd", x"3f2", x"3e7",
        x"3dd", x"3d2", x"3c7", x"3bc", x"3b2", x"3a7", x"39d", x"392",
        x"388", x"37d", x"373", x"369", x"35e", x"354", x"34a", x"340",
        x"336", x"32c", x"322", x"318", x"30e", x"304", x"2fa", x"2f0",
        x"2e7", x"2dd", x"2d3", x"2ca", x"2c0", x"2b7", x"2ad", x"2a4",
        x"29b", x"291", x"288", x"27f", x"276", x"26d", x"264", x"25b",
        x"252", x"249", x"241", x"238", x"22f", x"227", x"21e", x"216",
        x"20d", x"205", x"1fc", x"1f4", x"1ec", x"1e4", x"1dc", x"1d4",
        x"1cc", x"1c4", x"1bc", x"1b4", x"1ac", x"1a5", x"19d", x"196",
        x"18e", x"187", x"17f", x"178", x"171", x"16a", x"163", x"15b",
        x"154", x"14e", x"147", x"140", x"139", x"133", x"12c", x"125",
        x"11f", x"119", x"112", x"10c", x"106", x"100", x"0fa", x"0f4",
        x"0ee", x"0e8", x"0e2", x"0dc", x"0d7", x"0d1", x"0cc", x"0c6",
        x"0c1", x"0bc", x"0b6", x"0b1", x"0ac", x"0a7", x"0a2", x"09d",
        x"099", x"094", x"08f", x"08b", x"086", x"082", x"07d", x"079",
        x"075", x"071", x"06d", x"069", x"065", x"061", x"05d", x"059",
        x"056", x"052", x"04f", x"04b", x"048", x"045", x"041", x"03e",
        x"03b", x"038", x"035", x"033", x"030", x"02d", x"02b", x"028",
        x"026", x"023", x"021", x"01f", x"01d", x"01b", x"019", x"017",
        x"015", x"013", x"011", x"010", x"00e", x"00d", x"00b", x"00a",
        x"009", x"008", x"007", x"006", x"005", x"004", x"003", x"003",
        x"002", x"002", x"001", x"001", x"000", x"000", x"000", x"000",
        x"000", x"000", x"000", x"001", x"001", x"001", x"002", x"002",
        x"003", x"004", x"004", x"005", x"006", x"007", x"008", x"00a",
        x"00b", x"00c", x"00e", x"00f", x"011", x"012", x"014", x"016",
        x"018", x"01a", x"01c", x"01e", x"020", x"022", x"024", x"027",
        x"029", x"02c", x"02e", x"031", x"034", x"037", x"03a", x"03d",
        x"040", x"043", x"046", x"049", x"04d", x"050", x"054", x"057",
        x"05b", x"05f", x"063", x"067", x"06b", x"06f", x"073", x"077",
        x"07b", x"07f", x"084", x"088", x"08d", x"092", x"096", x"09b",
        x"0a0", x"0a5", x"0aa", x"0af", x"0b4", x"0b9", x"0be", x"0c4",
        x"0c9", x"0ce", x"0d4", x"0da", x"0df", x"0e5", x"0eb", x"0f1",
        x"0f7", x"0fd", x"103", x"109", x"10f", x"115", x"11c", x"122",
        x"129", x"12f", x"136", x"13d", x"143", x"14a", x"151", x"158",
        x"15f", x"166", x"16d", x"174", x"17c", x"183", x"18a", x"192",
        x"199", x"1a1", x"1a9", x"1b0", x"1b8", x"1c0", x"1c8", x"1d0",
        x"1d8", x"1e0", x"1e8", x"1f0", x"1f8", x"201", x"209", x"211",
        x"21a", x"222", x"22b", x"233", x"23c", x"245", x"24e", x"257",
        x"260", x"268", x"271", x"27b", x"284", x"28d", x"296", x"29f",
        x"2a9", x"2b2", x"2bc", x"2c5", x"2cf", x"2d8", x"2e2", x"2ec",
        x"2f5", x"2ff", x"309", x"313", x"31d", x"327", x"331", x"33b",
        x"345", x"34f", x"359", x"364", x"36e", x"378", x"383", x"38d",
        x"397", x"3a2", x"3ad", x"3b7", x"3c2", x"3cc", x"3d7", x"3e2",
        x"3ed", x"3f8", x"402", x"40d", x"418", x"423", x"42e", x"439",
        x"445", x"450", x"45b", x"466", x"471", x"47d", x"488", x"493",
        x"49f", x"4aa", x"4b6", x"4c1", x"4cd", x"4d8", x"4e4", x"4ef",
        x"4fb", x"507", x"512", x"51e", x"52a", x"535", x"541", x"54d",
        x"559", x"565", x"571", x"57d", x"589", x"595", x"5a1", x"5ad",
        x"5b9", x"5c5", x"5d1", x"5dd", x"5e9", x"5f5", x"601", x"60e",
        x"61a", x"626", x"632", x"63e", x"64b", x"657", x"663", x"670",
        x"67c", x"688", x"695", x"6a1", x"6ae", x"6ba", x"6c6", x"6d3",
        x"6df", x"6ec", x"6f8", x"705", x"711", x"71e", x"72a", x"737",
        x"743", x"750", x"75c", x"769", x"775", x"782", x"78e", x"79b",
        x"7a7", x"7b4", x"7c1", x"7cd", x"7da", x"7e6", x"7f3", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800",
        x"800", x"800", x"800", x"800", x"800", x"800", x"800", x"800"
    );
    signal tmp: std_logic_vector(11 downto 0);
begin

    ret: process (addr,clk) begin
        if (clk' event and clk = '1') then
            tmp <= ROM(conv_integer(addr));
        end if;
    end process;

    buff: process (tmp,en) begin
        if(en = '1') then
            data <= tmp;
        else
            data <= (others => 'Z');
        end if;
    end process buff;
end arch;
